magic
tech scmos
timestamp 1719641852
<< metal1 >>
rect 344 3603 346 3607
rect 350 3603 353 3607
rect 357 3603 360 3607
rect 1360 3603 1362 3607
rect 1366 3603 1369 3607
rect 1373 3603 1376 3607
rect 2384 3603 2386 3607
rect 2390 3603 2393 3607
rect 2397 3603 2400 3607
rect 3408 3603 3410 3607
rect 3414 3603 3417 3607
rect 3421 3603 3424 3607
rect 2450 3568 2451 3572
rect 3197 3568 3198 3572
rect 3310 3568 3321 3571
rect 2382 3558 2398 3561
rect 334 3548 369 3551
rect 550 3548 569 3551
rect 774 3548 809 3551
rect 1170 3548 1177 3551
rect 1402 3548 1417 3551
rect 1671 3548 1689 3551
rect 1895 3548 1929 3551
rect 2466 3548 2473 3551
rect 2866 3548 2873 3551
rect 2878 3548 2886 3551
rect 2926 3551 2929 3561
rect 3230 3561 3233 3568
rect 3318 3562 3321 3568
rect 2894 3548 2929 3551
rect 3214 3551 3217 3561
rect 3230 3558 3241 3561
rect 3202 3548 3217 3551
rect 3222 3548 3230 3551
rect 3270 3548 3289 3551
rect 3382 3548 3401 3551
rect 3406 3548 3422 3551
rect 3530 3548 3537 3551
rect 174 3538 177 3548
rect 2098 3538 2105 3541
rect 2394 3538 2417 3541
rect 2914 3538 2929 3541
rect 3142 3538 3158 3541
rect 3230 3538 3241 3541
rect 3278 3538 3286 3541
rect 3370 3538 3377 3541
rect 3518 3538 3529 3541
rect 2414 3528 2417 3538
rect 3518 3532 3521 3538
rect 3118 3528 3137 3531
rect 3154 3528 3166 3531
rect 3478 3521 3481 3528
rect 3478 3518 3489 3521
rect 848 3503 850 3507
rect 854 3503 857 3507
rect 861 3503 864 3507
rect 1880 3503 1882 3507
rect 1886 3503 1889 3507
rect 1893 3503 1896 3507
rect 2904 3503 2906 3507
rect 2910 3503 2913 3507
rect 2917 3503 2920 3507
rect 1334 3488 1350 3491
rect 2930 3488 2937 3491
rect 1694 3478 1710 3481
rect 2326 3478 2350 3481
rect 2190 3468 2206 3471
rect 2266 3468 2281 3471
rect 2814 3468 2825 3471
rect 2974 3468 2985 3471
rect 3006 3468 3014 3471
rect 3030 3468 3041 3471
rect 3166 3468 3185 3471
rect 222 3458 241 3461
rect 630 3452 633 3462
rect 1182 3458 1201 3461
rect 1242 3458 1254 3461
rect 1478 3458 1481 3468
rect 2286 3458 2313 3461
rect 2554 3458 2561 3461
rect 3010 3458 3025 3461
rect 3054 3458 3062 3461
rect 3070 3458 3078 3461
rect 3110 3458 3118 3461
rect 3302 3461 3305 3471
rect 3406 3471 3409 3481
rect 3406 3468 3438 3471
rect 3470 3468 3481 3471
rect 3302 3458 3310 3461
rect 3318 3458 3326 3461
rect 3390 3461 3393 3468
rect 3374 3458 3393 3461
rect 3478 3462 3481 3468
rect 3214 3448 3222 3451
rect 3498 3448 3505 3451
rect 3546 3448 3553 3451
rect 974 3438 982 3441
rect 3254 3438 3262 3441
rect 3366 3441 3370 3444
rect 3346 3438 3370 3441
rect 3194 3418 3195 3422
rect 3293 3418 3294 3422
rect 3397 3418 3398 3422
rect 344 3403 346 3407
rect 350 3403 353 3407
rect 357 3403 360 3407
rect 1360 3403 1362 3407
rect 1366 3403 1369 3407
rect 1373 3403 1376 3407
rect 2384 3403 2386 3407
rect 2390 3403 2393 3407
rect 2397 3403 2400 3407
rect 3408 3403 3410 3407
rect 3414 3403 3417 3407
rect 3421 3403 3424 3407
rect 298 3388 299 3392
rect 330 3388 331 3392
rect 378 3388 379 3392
rect 645 3388 646 3392
rect 674 3388 675 3392
rect 1274 3388 1275 3392
rect 2189 3388 2190 3392
rect 2954 3388 2955 3392
rect 934 3371 937 3381
rect 1302 3371 1305 3381
rect 934 3368 954 3371
rect 1286 3368 1305 3371
rect 1590 3368 1601 3371
rect 2774 3368 2782 3371
rect 3218 3368 3241 3371
rect 3286 3368 3297 3371
rect 3434 3368 3449 3371
rect 3746 3368 3769 3371
rect 1590 3362 1593 3368
rect 1606 3366 1610 3368
rect 3294 3362 3297 3368
rect 686 3358 705 3361
rect 1978 3358 1985 3361
rect 3174 3352 3177 3361
rect 3326 3358 3337 3361
rect 46 3348 54 3351
rect 290 3348 297 3351
rect 322 3348 329 3351
rect 650 3348 673 3351
rect 966 3348 993 3351
rect 1046 3348 1054 3351
rect 1078 3348 1086 3351
rect 1358 3348 1366 3351
rect 3158 3348 3174 3351
rect 3386 3348 3393 3351
rect 3470 3348 3489 3351
rect 3518 3348 3529 3351
rect 658 3338 665 3341
rect 986 3338 993 3341
rect 1326 3341 1329 3348
rect 3486 3342 3489 3348
rect 3526 3342 3529 3348
rect 1326 3338 1345 3341
rect 1682 3338 1689 3341
rect 1774 3338 1782 3341
rect 2914 3338 2929 3341
rect 2974 3338 2993 3341
rect 2998 3338 3009 3341
rect 3502 3338 3510 3341
rect 2998 3332 3001 3338
rect 62 3328 70 3331
rect 2430 3328 2438 3331
rect 3270 3331 3273 3338
rect 3262 3328 3273 3331
rect 3490 3328 3497 3331
rect 3502 3328 3505 3338
rect 3702 3328 3710 3331
rect 3758 3331 3761 3338
rect 3758 3328 3769 3331
rect 2394 3318 2395 3322
rect 2418 3318 2425 3321
rect 3058 3318 3060 3322
rect 3098 3318 3100 3322
rect 3181 3318 3182 3322
rect 848 3303 850 3307
rect 854 3303 857 3307
rect 861 3303 864 3307
rect 1880 3303 1882 3307
rect 1886 3303 1889 3307
rect 1893 3303 1896 3307
rect 2904 3303 2906 3307
rect 2910 3303 2913 3307
rect 2917 3303 2920 3307
rect 418 3288 433 3291
rect 1366 3288 1374 3291
rect 2900 3288 2902 3292
rect 2342 3278 2350 3281
rect 2386 3278 2398 3281
rect 2994 3278 3001 3281
rect 3754 3278 3761 3281
rect 482 3268 489 3271
rect 646 3268 654 3271
rect 1454 3268 1473 3271
rect 1598 3268 1606 3271
rect 1638 3268 1649 3271
rect 1674 3268 1681 3271
rect 2438 3268 2446 3271
rect 2454 3268 2473 3271
rect 2534 3268 2545 3271
rect 2582 3268 2601 3271
rect 3078 3268 3086 3271
rect 3134 3268 3153 3271
rect 3226 3268 3233 3271
rect 3298 3268 3305 3271
rect 1638 3262 1641 3268
rect 3366 3268 3393 3271
rect 3398 3268 3406 3271
rect 3690 3268 3697 3271
rect 22 3258 41 3261
rect 474 3258 497 3261
rect 542 3258 561 3261
rect 566 3258 593 3261
rect 618 3258 625 3261
rect 822 3258 830 3261
rect 1014 3258 1018 3262
rect 1242 3258 1249 3261
rect 1438 3258 1457 3261
rect 2286 3258 2294 3261
rect 2354 3258 2361 3261
rect 2462 3258 2470 3261
rect 2558 3258 2566 3261
rect 2602 3258 2609 3261
rect 2658 3258 2665 3261
rect 3254 3258 3273 3261
rect 3462 3258 3470 3261
rect 3682 3258 3705 3261
rect 734 3248 745 3251
rect 1014 3252 1017 3258
rect 1542 3252 1546 3254
rect 1310 3248 1329 3251
rect 2282 3248 2286 3252
rect 3182 3251 3185 3258
rect 3182 3248 3193 3251
rect 3242 3248 3246 3252
rect 3254 3248 3257 3258
rect 3402 3248 3425 3251
rect 526 3238 534 3241
rect 3126 3241 3129 3248
rect 3606 3246 3610 3248
rect 1406 3238 1426 3241
rect 3126 3238 3137 3241
rect 3606 3238 3614 3241
rect 722 3228 723 3232
rect 1262 3228 1265 3238
rect 1406 3228 1409 3238
rect 3162 3218 3163 3222
rect 3490 3218 3491 3222
rect 3677 3218 3678 3222
rect 344 3203 346 3207
rect 350 3203 353 3207
rect 357 3203 360 3207
rect 1360 3203 1362 3207
rect 1366 3203 1369 3207
rect 1373 3203 1376 3207
rect 2384 3203 2386 3207
rect 2390 3203 2393 3207
rect 2397 3203 2400 3207
rect 3408 3203 3410 3207
rect 3414 3203 3417 3207
rect 3421 3203 3424 3207
rect 773 3188 774 3192
rect 2037 3188 2038 3192
rect 2178 3188 2179 3192
rect 2293 3188 2294 3192
rect 2650 3188 2651 3192
rect 738 3168 750 3171
rect 878 3171 881 3181
rect 846 3168 881 3171
rect 1358 3168 1382 3171
rect 1446 3171 1449 3181
rect 1430 3168 1449 3171
rect 1798 3168 1809 3171
rect 2213 3168 2214 3172
rect 2330 3168 2337 3171
rect 2390 3168 2398 3171
rect 3266 3168 3267 3172
rect 3702 3168 3718 3171
rect 918 3166 922 3168
rect 718 3158 729 3161
rect 986 3158 990 3162
rect 1518 3161 1521 3168
rect 1542 3166 1546 3168
rect 1798 3162 1801 3168
rect 1814 3166 1818 3168
rect 3702 3166 3706 3168
rect 1518 3158 1537 3161
rect 918 3148 929 3151
rect 970 3148 977 3151
rect 918 3142 921 3148
rect 1126 3142 1129 3151
rect 1398 3148 1414 3151
rect 1422 3148 1430 3151
rect 1486 3148 1494 3151
rect 1678 3148 1686 3151
rect 1742 3151 1746 3154
rect 1742 3148 1761 3151
rect 1870 3151 1873 3161
rect 1878 3158 1913 3161
rect 1854 3148 1873 3151
rect 1890 3148 1921 3151
rect 1966 3151 1969 3161
rect 1950 3148 1969 3151
rect 1986 3148 2009 3151
rect 2082 3148 2089 3151
rect 2094 3148 2102 3151
rect 2150 3148 2177 3151
rect 2278 3151 2281 3161
rect 2418 3158 2425 3161
rect 2262 3148 2281 3151
rect 2402 3148 2433 3151
rect 2490 3148 2497 3151
rect 2502 3148 2510 3151
rect 2578 3148 2585 3151
rect 2590 3148 2617 3151
rect 2662 3151 2665 3161
rect 3122 3158 3126 3162
rect 2662 3148 2681 3151
rect 2894 3148 2918 3151
rect 2938 3148 2945 3151
rect 2974 3148 2998 3151
rect 3006 3148 3017 3151
rect 3074 3148 3081 3151
rect 3126 3148 3134 3151
rect 3198 3148 3217 3151
rect 3350 3151 3353 3161
rect 3382 3158 3390 3161
rect 3414 3158 3438 3161
rect 3322 3148 3353 3151
rect 3366 3148 3374 3151
rect 3494 3148 3513 3151
rect 946 3138 953 3141
rect 1690 3138 1697 3141
rect 1830 3138 1838 3141
rect 2102 3138 2110 3141
rect 2478 3138 2489 3141
rect 2526 3138 2545 3141
rect 2942 3138 2945 3148
rect 3014 3142 3017 3148
rect 2994 3138 3001 3141
rect 3070 3138 3078 3141
rect 3142 3141 3145 3148
rect 3134 3138 3145 3141
rect 3170 3138 3177 3141
rect 3198 3138 3201 3148
rect 3406 3138 3414 3141
rect 3606 3138 3633 3141
rect 1358 3128 1393 3131
rect 2854 3128 2862 3131
rect 914 3118 915 3122
rect 2117 3118 2118 3122
rect 2237 3118 2238 3122
rect 3550 3118 3558 3121
rect 848 3103 850 3107
rect 854 3103 857 3107
rect 861 3103 864 3107
rect 1880 3103 1882 3107
rect 1886 3103 1889 3107
rect 1893 3103 1896 3107
rect 2904 3103 2906 3107
rect 2910 3103 2913 3107
rect 2917 3103 2920 3107
rect 1717 3088 1718 3092
rect 2194 3088 2195 3092
rect 2602 3088 2603 3092
rect 206 3072 209 3081
rect 1134 3072 1137 3081
rect 1498 3078 1513 3081
rect 2002 3078 2009 3081
rect 2638 3078 2649 3081
rect 214 3068 222 3071
rect 458 3068 465 3071
rect 486 3062 489 3071
rect 706 3068 721 3071
rect 1150 3068 1158 3071
rect 1654 3068 1662 3071
rect 1686 3068 1694 3071
rect 2018 3068 2025 3071
rect 2066 3068 2073 3071
rect 682 3058 689 3061
rect 842 3058 849 3061
rect 1466 3058 1473 3061
rect 1726 3058 1734 3061
rect 2026 3058 2033 3061
rect 2126 3061 2129 3071
rect 2126 3058 2134 3061
rect 2158 3061 2161 3071
rect 2270 3062 2273 3071
rect 2978 3068 2985 3071
rect 3158 3068 3169 3071
rect 3190 3068 3201 3071
rect 3218 3068 3225 3071
rect 3294 3062 3297 3071
rect 3342 3068 3361 3071
rect 3410 3068 3425 3071
rect 3630 3068 3638 3071
rect 2158 3058 2185 3061
rect 2230 3058 2238 3061
rect 2322 3058 2329 3061
rect 2518 3058 2545 3061
rect 2558 3058 2577 3061
rect 2706 3058 2713 3061
rect 3306 3058 3313 3061
rect 3490 3058 3497 3061
rect 3514 3058 3521 3061
rect 242 3048 246 3052
rect 2182 3052 2185 3058
rect 1354 3048 1377 3051
rect 1750 3048 1758 3051
rect 1774 3048 1782 3051
rect 2458 3048 2462 3052
rect 2558 3048 2561 3058
rect 3466 3048 3470 3052
rect 3694 3051 3697 3058
rect 3594 3048 3609 3051
rect 3694 3048 3705 3051
rect 1134 3041 1137 3048
rect 1134 3038 1145 3041
rect 2710 3038 2718 3041
rect 3522 3038 3523 3042
rect 2546 3028 2547 3032
rect 3066 3018 3067 3022
rect 3253 3018 3254 3022
rect 3314 3018 3315 3022
rect 3621 3018 3622 3022
rect 3682 3018 3683 3022
rect 3757 3018 3758 3022
rect 344 3003 346 3007
rect 350 3003 353 3007
rect 357 3003 360 3007
rect 1360 3003 1362 3007
rect 1366 3003 1369 3007
rect 1373 3003 1376 3007
rect 2384 3003 2386 3007
rect 2390 3003 2393 3007
rect 2397 3003 2400 3007
rect 3408 3003 3410 3007
rect 3414 3003 3417 3007
rect 3421 3003 3424 3007
rect 525 2988 526 2992
rect 2125 2988 2126 2992
rect 2398 2988 2414 2991
rect 2466 2988 2467 2992
rect 2202 2978 2203 2982
rect 3342 2972 3345 2981
rect 1322 2968 1323 2972
rect 1358 2968 1366 2971
rect 894 2966 898 2968
rect 966 2966 970 2968
rect 974 2958 982 2961
rect 1230 2961 1233 2968
rect 1358 2966 1362 2968
rect 1230 2958 1241 2961
rect 1334 2958 1353 2961
rect 1626 2958 1633 2961
rect 822 2951 826 2954
rect 822 2948 841 2951
rect 926 2951 930 2954
rect 926 2948 945 2951
rect 1598 2951 1602 2954
rect 1694 2951 1697 2958
rect 2154 2958 2158 2962
rect 2434 2958 2438 2962
rect 1598 2948 1617 2951
rect 1686 2948 1697 2951
rect 2014 2948 2022 2951
rect 2038 2948 2054 2951
rect 2074 2948 2081 2951
rect 2186 2948 2201 2951
rect 2238 2948 2246 2951
rect 2358 2948 2374 2951
rect 2458 2948 2465 2951
rect 2486 2951 2489 2961
rect 2494 2958 2513 2961
rect 2482 2948 2489 2951
rect 2514 2948 2521 2951
rect 2526 2948 2553 2951
rect 2926 2948 2929 2958
rect 3334 2961 3338 2964
rect 3334 2958 3342 2961
rect 3430 2958 3441 2961
rect 3500 2958 3502 2962
rect 3738 2958 3745 2961
rect 3310 2948 3321 2951
rect 3430 2951 3433 2958
rect 3406 2948 3433 2951
rect 3534 2948 3545 2951
rect 578 2938 585 2941
rect 854 2938 862 2941
rect 874 2938 881 2941
rect 1622 2938 1630 2941
rect 2018 2938 2025 2941
rect 2166 2938 2177 2941
rect 2222 2941 2225 2948
rect 3318 2942 3321 2948
rect 3542 2942 3545 2948
rect 2222 2938 2233 2941
rect 2242 2938 2249 2941
rect 2274 2938 2281 2941
rect 2298 2938 2321 2941
rect 2334 2938 2350 2941
rect 3598 2938 3625 2941
rect 1230 2928 1233 2938
rect 2758 2928 2766 2931
rect 890 2918 891 2922
rect 1370 2918 1385 2921
rect 1637 2918 1638 2922
rect 2061 2918 2062 2922
rect 2258 2918 2259 2922
rect 2282 2918 2283 2922
rect 3141 2918 3142 2922
rect 3165 2918 3166 2922
rect 3212 2918 3214 2922
rect 3666 2918 3673 2921
rect 848 2903 850 2907
rect 854 2903 857 2907
rect 861 2903 864 2907
rect 1880 2903 1882 2907
rect 1886 2903 1889 2907
rect 1893 2903 1896 2907
rect 2904 2903 2906 2907
rect 2910 2903 2913 2907
rect 2917 2903 2920 2907
rect 882 2888 889 2891
rect 1466 2888 1473 2891
rect 2490 2888 2491 2892
rect 3458 2888 3459 2892
rect 1494 2872 1497 2881
rect 630 2868 641 2871
rect 734 2868 742 2871
rect 1286 2868 1294 2871
rect 1354 2868 1361 2871
rect 2006 2868 2014 2871
rect 2130 2868 2137 2871
rect 2230 2868 2241 2871
rect 2410 2868 2433 2871
rect 2526 2868 2537 2871
rect 226 2858 233 2861
rect 374 2858 377 2868
rect 686 2858 694 2861
rect 1074 2858 1081 2861
rect 1374 2858 1382 2861
rect 1422 2858 1425 2868
rect 1446 2858 1449 2868
rect 2230 2862 2233 2868
rect 1726 2858 1734 2861
rect 1986 2858 1993 2861
rect 2030 2858 2049 2861
rect 2086 2858 2102 2861
rect 2170 2858 2177 2861
rect 2182 2858 2209 2861
rect 2358 2858 2385 2861
rect 2494 2858 2513 2861
rect 2574 2861 2577 2871
rect 2626 2868 2633 2871
rect 2750 2871 2753 2881
rect 2994 2878 3009 2881
rect 3426 2878 3433 2881
rect 2734 2868 2753 2871
rect 2778 2868 2785 2871
rect 3438 2868 3449 2871
rect 3658 2868 3665 2871
rect 3734 2868 3753 2871
rect 2574 2858 2590 2861
rect 3154 2858 3169 2861
rect 3286 2858 3297 2861
rect 3598 2858 3617 2861
rect 3630 2858 3649 2861
rect 3686 2858 3705 2861
rect 3710 2858 3737 2861
rect 3750 2858 3753 2868
rect 66 2848 70 2852
rect 130 2848 134 2852
rect 694 2848 705 2851
rect 1058 2848 1065 2851
rect 2046 2848 2049 2858
rect 2494 2848 2497 2858
rect 3614 2848 3617 2858
rect 3686 2848 3689 2858
rect 414 2838 430 2841
rect 786 2838 787 2842
rect 1270 2841 1273 2848
rect 1054 2838 1074 2841
rect 1270 2838 1281 2841
rect 1326 2838 1342 2841
rect 3002 2838 3017 2841
rect 3438 2838 3446 2841
rect 3594 2838 3595 2842
rect 1054 2828 1057 2838
rect 3236 2828 3238 2832
rect 3365 2828 3366 2832
rect 853 2818 854 2822
rect 2277 2818 2278 2822
rect 3130 2818 3131 2822
rect 3394 2818 3395 2822
rect 3500 2818 3502 2822
rect 344 2803 346 2807
rect 350 2803 353 2807
rect 357 2803 360 2807
rect 1360 2803 1362 2807
rect 1366 2803 1369 2807
rect 1373 2803 1376 2807
rect 2384 2803 2386 2807
rect 2390 2803 2393 2807
rect 2397 2803 2400 2807
rect 3408 2803 3410 2807
rect 3414 2803 3417 2807
rect 3421 2803 3424 2807
rect 682 2788 683 2792
rect 746 2788 747 2792
rect 1845 2788 1846 2792
rect 2818 2788 2819 2792
rect 650 2778 651 2782
rect 598 2768 606 2771
rect 710 2771 713 2781
rect 925 2778 926 2782
rect 694 2768 713 2771
rect 802 2768 817 2771
rect 1994 2768 1995 2772
rect 3702 2771 3705 2781
rect 3686 2768 3705 2771
rect 942 2766 946 2768
rect 842 2758 846 2762
rect 854 2758 862 2761
rect 1002 2758 1006 2762
rect 22 2748 41 2751
rect 630 2748 649 2751
rect 982 2748 990 2751
rect 1370 2748 1377 2751
rect 1502 2748 1510 2751
rect 1750 2751 1754 2754
rect 1830 2751 1833 2761
rect 2786 2758 2790 2762
rect 1750 2748 1769 2751
rect 1814 2748 1833 2751
rect 1886 2748 1910 2751
rect 1926 2748 1934 2751
rect 2266 2748 2273 2751
rect 2278 2748 2286 2751
rect 2326 2748 2353 2751
rect 2390 2748 2414 2751
rect 2446 2748 2454 2751
rect 2802 2748 2817 2751
rect 2894 2748 2910 2751
rect 3078 2748 3081 2758
rect 3274 2748 3281 2751
rect 3506 2748 3513 2751
rect 3570 2748 3577 2751
rect 3758 2748 3769 2751
rect 622 2738 625 2748
rect 942 2741 945 2748
rect 942 2738 953 2741
rect 1390 2738 1398 2741
rect 1854 2738 1873 2741
rect 1898 2738 1913 2741
rect 1934 2738 1953 2741
rect 1974 2738 1985 2741
rect 2054 2738 2070 2741
rect 2702 2738 2713 2741
rect 2734 2738 2753 2741
rect 2874 2738 2881 2741
rect 3262 2741 3265 2748
rect 3758 2742 3761 2748
rect 3255 2738 3265 2741
rect 3350 2738 3369 2741
rect 3646 2738 3662 2741
rect 1962 2728 1969 2731
rect 3470 2728 3481 2731
rect 1341 2718 1342 2722
rect 1789 2718 1790 2722
rect 3332 2718 3334 2722
rect 848 2703 850 2707
rect 854 2703 857 2707
rect 861 2703 864 2707
rect 1880 2703 1882 2707
rect 1886 2703 1889 2707
rect 1893 2703 1896 2707
rect 2904 2703 2906 2707
rect 2910 2703 2913 2707
rect 2917 2703 2920 2707
rect 853 2688 854 2692
rect 1542 2678 1561 2681
rect 2654 2678 2673 2681
rect 2710 2678 2729 2681
rect 2878 2678 2897 2681
rect 6 2662 9 2671
rect 322 2668 329 2671
rect 346 2668 361 2671
rect 406 2662 409 2671
rect 606 2668 614 2671
rect 654 2668 670 2671
rect 734 2668 742 2671
rect 1487 2668 1505 2671
rect 1598 2668 1609 2671
rect 1886 2668 1902 2671
rect 2122 2668 2129 2671
rect 2374 2668 2382 2671
rect 2394 2668 2401 2671
rect 2814 2662 2817 2671
rect 2870 2668 2878 2671
rect 3298 2668 3305 2671
rect 3358 2668 3377 2671
rect 3454 2668 3470 2671
rect 3490 2668 3497 2671
rect 3718 2668 3729 2671
rect 334 2658 350 2661
rect 1022 2658 1030 2661
rect 721 2648 726 2652
rect 937 2648 942 2652
rect 1334 2652 1337 2661
rect 1854 2658 1873 2661
rect 2086 2658 2094 2661
rect 2270 2658 2289 2661
rect 2302 2658 2329 2661
rect 2334 2658 2361 2661
rect 2378 2658 2409 2661
rect 2414 2658 2422 2661
rect 2750 2658 2758 2661
rect 2906 2658 2937 2661
rect 3262 2658 3265 2668
rect 3318 2658 3326 2661
rect 3342 2658 3350 2661
rect 3478 2658 3505 2661
rect 3634 2658 3649 2661
rect 3654 2658 3662 2661
rect 3678 2658 3689 2661
rect 3694 2658 3702 2661
rect 1854 2648 1857 2658
rect 2286 2648 2289 2658
rect 3550 2648 3558 2651
rect 3622 2648 3630 2651
rect 3750 2648 3774 2651
rect 846 2642 850 2644
rect 1110 2641 1114 2644
rect 1102 2638 1114 2641
rect 2773 2638 2774 2642
rect 3538 2638 3577 2641
rect 2301 2628 2302 2632
rect 2154 2618 2155 2622
rect 3157 2618 3158 2622
rect 3221 2618 3222 2622
rect 3386 2618 3387 2622
rect 3422 2618 3438 2621
rect 3506 2618 3507 2622
rect 3738 2618 3739 2622
rect 344 2603 346 2607
rect 350 2603 353 2607
rect 357 2603 360 2607
rect 1360 2603 1362 2607
rect 1366 2603 1369 2607
rect 1373 2603 1376 2607
rect 2384 2603 2386 2607
rect 2390 2603 2393 2607
rect 2397 2603 2400 2607
rect 3408 2603 3410 2607
rect 3414 2603 3417 2607
rect 3421 2603 3424 2607
rect 1221 2588 1222 2592
rect 2426 2588 2427 2592
rect 2746 2588 2747 2592
rect 2810 2588 2811 2592
rect 2877 2588 2878 2592
rect 2938 2588 2939 2592
rect 2381 2578 2382 2582
rect 2586 2578 2587 2582
rect 2717 2568 2718 2572
rect 794 2558 798 2562
rect 1078 2552 1081 2561
rect 1514 2558 1521 2561
rect 2554 2558 2558 2562
rect 2650 2558 2654 2562
rect 2758 2558 2769 2561
rect 22 2548 41 2551
rect 590 2548 617 2551
rect 878 2548 886 2551
rect 950 2548 958 2551
rect 1058 2548 1073 2551
rect 1902 2548 1910 2551
rect 2462 2548 2489 2551
rect 2494 2548 2502 2551
rect 2546 2548 2553 2551
rect 2578 2548 2585 2551
rect 2622 2548 2638 2551
rect 2674 2548 2681 2551
rect 2834 2548 2841 2551
rect 2846 2548 2862 2551
rect 2950 2551 2953 2561
rect 3762 2558 3766 2562
rect 2914 2548 2937 2551
rect 2950 2548 2969 2551
rect 3010 2548 3017 2551
rect 574 2538 577 2548
rect 1479 2538 1494 2541
rect 1510 2538 1513 2548
rect 3062 2542 3065 2551
rect 3150 2548 3158 2551
rect 3206 2548 3225 2551
rect 3246 2548 3265 2551
rect 3378 2548 3385 2551
rect 3422 2548 3446 2551
rect 3606 2548 3614 2551
rect 3630 2548 3638 2551
rect 3674 2548 3681 2551
rect 1790 2538 1798 2541
rect 1854 2538 1889 2541
rect 2410 2538 2417 2541
rect 3002 2538 3009 2541
rect 3102 2538 3129 2541
rect 3142 2538 3169 2541
rect 3178 2538 3185 2541
rect 3266 2538 3273 2541
rect 3298 2538 3305 2541
rect 3358 2538 3377 2541
rect 3454 2538 3473 2541
rect 3546 2538 3561 2541
rect 1726 2528 1734 2531
rect 1738 2528 1745 2531
rect 1750 2528 1758 2531
rect 3282 2528 3286 2532
rect 3346 2528 3353 2531
rect 1074 2518 1075 2522
rect 1285 2518 1286 2522
rect 2117 2518 2118 2522
rect 3141 2518 3142 2522
rect 3653 2518 3654 2522
rect 848 2503 850 2507
rect 854 2503 857 2507
rect 861 2503 864 2507
rect 1880 2503 1882 2507
rect 1886 2503 1889 2507
rect 1893 2503 1896 2507
rect 2904 2503 2906 2507
rect 2910 2503 2913 2507
rect 2917 2503 2920 2507
rect 1014 2478 1030 2481
rect 2470 2478 2481 2481
rect 1014 2472 1017 2478
rect 678 2462 681 2471
rect 722 2468 729 2471
rect 1246 2468 1265 2471
rect 1734 2471 1737 2478
rect 1734 2468 1745 2471
rect 1806 2468 1825 2471
rect 1898 2468 1905 2471
rect 2142 2468 2150 2471
rect 2314 2468 2329 2471
rect 2766 2468 2790 2471
rect 2818 2468 2825 2471
rect 3006 2468 3014 2471
rect 3242 2468 3249 2471
rect 3318 2468 3337 2471
rect 3402 2468 3409 2471
rect 3418 2468 3441 2471
rect 58 2458 65 2461
rect 742 2458 750 2461
rect 794 2458 801 2461
rect 818 2458 825 2461
rect 1042 2458 1049 2461
rect 1074 2458 1081 2461
rect 1146 2458 1153 2461
rect 1782 2458 1793 2461
rect 1838 2458 1846 2461
rect 1858 2458 1865 2461
rect 1918 2458 1937 2461
rect 1974 2458 1993 2461
rect 2278 2458 2297 2461
rect 2302 2458 2318 2461
rect 2390 2461 2393 2468
rect 2390 2458 2417 2461
rect 2438 2458 2454 2461
rect 66 2448 70 2452
rect 750 2448 761 2451
rect 1878 2448 1913 2451
rect 1918 2448 1921 2458
rect 1990 2448 1993 2458
rect 1998 2448 2017 2451
rect 2082 2448 2086 2452
rect 2094 2448 2113 2451
rect 2750 2448 2758 2451
rect 3554 2448 3561 2451
rect 790 2442 794 2444
rect 642 2438 665 2441
rect 1022 2441 1026 2444
rect 1014 2438 1026 2441
rect 1198 2438 1206 2441
rect 1698 2438 1699 2442
rect 917 2428 918 2432
rect 3450 2428 3451 2432
rect 3732 2418 3734 2422
rect 344 2403 346 2407
rect 350 2403 353 2407
rect 357 2403 360 2407
rect 1360 2403 1362 2407
rect 1366 2403 1369 2407
rect 1373 2403 1376 2407
rect 2384 2403 2386 2407
rect 2390 2403 2393 2407
rect 2397 2403 2400 2407
rect 3408 2403 3410 2407
rect 3414 2403 3417 2407
rect 3421 2403 3424 2407
rect 498 2388 499 2392
rect 986 2388 987 2392
rect 1258 2388 1259 2392
rect 2050 2388 2051 2392
rect 2754 2388 2755 2392
rect 530 2368 531 2372
rect 690 2368 691 2372
rect 750 2371 753 2381
rect 734 2368 753 2371
rect 3446 2371 3449 2381
rect 3674 2378 3675 2382
rect 3446 2368 3481 2371
rect 3734 2368 3742 2371
rect 1562 2358 1566 2362
rect 46 2348 65 2351
rect 490 2348 497 2351
rect 558 2348 577 2351
rect 802 2348 809 2351
rect 814 2348 822 2351
rect 1022 2348 1030 2351
rect 1238 2348 1257 2351
rect 1614 2351 1617 2361
rect 1622 2358 1641 2361
rect 2666 2358 2670 2362
rect 2678 2352 2681 2361
rect 2766 2358 2777 2361
rect 3094 2358 3105 2361
rect 1598 2348 1617 2351
rect 1858 2348 1865 2351
rect 1890 2348 1897 2351
rect 1946 2348 1961 2351
rect 2022 2348 2030 2351
rect 2042 2348 2049 2351
rect 2614 2348 2625 2351
rect 2722 2348 2729 2351
rect 391 2338 425 2341
rect 1334 2341 1337 2348
rect 1334 2338 1345 2341
rect 1670 2341 1673 2348
rect 1670 2338 1681 2341
rect 1710 2338 1718 2341
rect 1910 2338 1929 2341
rect 2738 2338 2745 2341
rect 2850 2338 2857 2341
rect 2874 2338 2905 2341
rect 3166 2338 3174 2341
rect 3210 2338 3217 2341
rect 3234 2338 3249 2341
rect 3266 2338 3281 2341
rect 3290 2338 3313 2341
rect 3366 2338 3385 2341
rect 3502 2338 3521 2341
rect 3558 2338 3577 2341
rect 3646 2338 3665 2341
rect 790 2332 793 2338
rect 786 2328 793 2332
rect 1350 2328 1374 2331
rect 1874 2328 1897 2331
rect 2574 2328 2593 2331
rect 2710 2328 2718 2331
rect 2830 2328 2849 2331
rect 3194 2328 3198 2332
rect 1037 2318 1038 2322
rect 3406 2318 3414 2321
rect 3484 2318 3486 2322
rect 848 2303 850 2307
rect 854 2303 857 2307
rect 861 2303 864 2307
rect 1880 2303 1882 2307
rect 1886 2303 1889 2307
rect 1893 2303 1896 2307
rect 2904 2303 2906 2307
rect 2910 2303 2913 2307
rect 2917 2303 2920 2307
rect 1194 2288 1201 2291
rect 1466 2288 1467 2292
rect 2386 2288 2401 2291
rect 3226 2288 3227 2292
rect 1174 2272 1177 2281
rect 2518 2278 2529 2281
rect 2826 2278 2833 2281
rect 206 2268 217 2271
rect 426 2268 433 2271
rect 926 2268 945 2271
rect 1038 2268 1057 2271
rect 206 2262 209 2268
rect 1422 2262 1425 2271
rect 94 2258 102 2261
rect 230 2258 238 2261
rect 438 2258 457 2261
rect 638 2258 642 2262
rect 1006 2258 1025 2261
rect 1082 2258 1089 2261
rect 1438 2258 1446 2261
rect 1454 2261 1457 2271
rect 1726 2268 1734 2271
rect 1870 2268 1881 2271
rect 1906 2268 1913 2271
rect 1990 2268 2009 2271
rect 2086 2268 2097 2271
rect 2178 2268 2185 2271
rect 1870 2262 1873 2268
rect 2094 2262 2097 2268
rect 2486 2262 2489 2271
rect 2834 2268 2841 2271
rect 3046 2268 3054 2271
rect 3154 2268 3161 2271
rect 3238 2268 3265 2271
rect 3294 2268 3302 2271
rect 3306 2268 3321 2271
rect 3350 2268 3358 2271
rect 3374 2268 3393 2271
rect 3446 2268 3454 2271
rect 1450 2258 1457 2261
rect 1470 2258 1489 2261
rect 1718 2258 1745 2261
rect 1806 2258 1833 2261
rect 2066 2258 2073 2261
rect 2550 2261 2553 2268
rect 2550 2258 2561 2261
rect 2626 2258 2633 2261
rect 2846 2258 2854 2261
rect 3026 2258 3038 2261
rect 3102 2258 3110 2261
rect 3182 2258 3201 2261
rect 3382 2258 3390 2261
rect 3490 2258 3497 2261
rect 3502 2258 3518 2261
rect 114 2248 118 2252
rect 638 2252 641 2258
rect 1022 2248 1025 2258
rect 1470 2248 1473 2258
rect 1770 2248 1774 2252
rect 3078 2248 3089 2251
rect 3098 2248 3102 2252
rect 3414 2248 3430 2251
rect 2445 2238 2446 2242
rect 2914 2218 2929 2221
rect 3402 2218 3403 2222
rect 3706 2218 3707 2222
rect 344 2203 346 2207
rect 350 2203 353 2207
rect 357 2203 360 2207
rect 1360 2203 1362 2207
rect 1366 2203 1369 2207
rect 1373 2203 1376 2207
rect 2384 2203 2386 2207
rect 2390 2203 2393 2207
rect 2397 2203 2400 2207
rect 3408 2203 3410 2207
rect 3414 2203 3417 2207
rect 3421 2203 3424 2207
rect 757 2188 758 2192
rect 1386 2188 1401 2191
rect 1530 2188 1531 2192
rect 2293 2188 2294 2192
rect 2466 2188 2467 2192
rect 2498 2188 2499 2192
rect 2562 2188 2563 2192
rect 3514 2188 3515 2192
rect 3546 2188 3547 2192
rect 3698 2188 3699 2192
rect 726 2171 729 2181
rect 726 2168 746 2171
rect 790 2171 793 2181
rect 790 2168 810 2171
rect 1638 2168 1649 2171
rect 1646 2162 1649 2168
rect 530 2158 534 2162
rect 542 2158 553 2161
rect 1158 2158 1177 2161
rect 22 2148 30 2151
rect 510 2148 529 2151
rect 670 2148 678 2151
rect 1170 2148 1185 2151
rect 1494 2151 1497 2158
rect 1542 2151 1545 2161
rect 1486 2148 1497 2151
rect 1502 2148 1529 2151
rect 1542 2148 1561 2151
rect 1614 2148 1630 2151
rect 1670 2151 1673 2161
rect 1654 2148 1673 2151
rect 1686 2148 1713 2151
rect 1718 2148 1745 2151
rect 1750 2148 1758 2151
rect 1830 2151 1833 2161
rect 1922 2158 1926 2162
rect 1954 2158 1958 2162
rect 2386 2158 2390 2162
rect 2714 2158 2718 2162
rect 1814 2148 1833 2151
rect 1886 2148 1913 2151
rect 1978 2148 1985 2151
rect 2334 2148 2342 2151
rect 2402 2148 2433 2151
rect 2598 2148 2606 2151
rect 2654 2148 2662 2151
rect 2730 2148 2745 2151
rect 2814 2151 2817 2161
rect 2798 2148 2817 2151
rect 3190 2148 3209 2151
rect 3294 2148 3305 2151
rect 3450 2148 3457 2151
rect 3462 2148 3470 2151
rect 466 2138 481 2141
rect 1126 2138 1129 2148
rect 1910 2142 1913 2148
rect 3294 2142 3297 2148
rect 1478 2138 1486 2141
rect 1574 2138 1601 2141
rect 1758 2138 1766 2141
rect 1854 2138 1873 2141
rect 2398 2138 2414 2141
rect 2542 2138 2550 2141
rect 3154 2138 3169 2141
rect 3250 2138 3265 2141
rect 3338 2138 3361 2141
rect 3486 2138 3505 2141
rect 502 2128 505 2138
rect 3178 2128 3182 2132
rect 1477 2118 1478 2122
rect 3740 2118 3742 2122
rect 848 2103 850 2107
rect 854 2103 857 2107
rect 861 2103 864 2107
rect 1880 2103 1882 2107
rect 1886 2103 1889 2107
rect 1893 2103 1896 2107
rect 2904 2103 2906 2107
rect 2910 2103 2913 2107
rect 2917 2103 2920 2107
rect 1196 2088 1198 2092
rect 3277 2088 3278 2092
rect 3597 2088 3598 2092
rect 3682 2088 3689 2091
rect 1242 2078 1249 2081
rect 606 2068 617 2071
rect 1230 2068 1246 2071
rect 1430 2068 1441 2071
rect 1462 2062 1465 2071
rect 1526 2071 1529 2081
rect 1906 2078 1913 2081
rect 2358 2078 2377 2081
rect 2630 2078 2641 2081
rect 2942 2078 2953 2081
rect 2998 2078 3009 2081
rect 3574 2081 3577 2088
rect 3566 2078 3577 2081
rect 2950 2072 2953 2078
rect 1526 2068 1545 2071
rect 1730 2068 1737 2071
rect 1934 2068 1953 2071
rect 46 2058 54 2061
rect 494 2058 510 2061
rect 662 2058 670 2061
rect 886 2058 894 2061
rect 1470 2058 1473 2068
rect 1934 2062 1937 2068
rect 1798 2058 1817 2061
rect 2158 2061 2161 2071
rect 2330 2068 2337 2071
rect 2418 2068 2425 2071
rect 2570 2068 2577 2071
rect 2903 2068 2937 2071
rect 3054 2071 3057 2078
rect 3054 2068 3073 2071
rect 3110 2068 3118 2071
rect 3286 2068 3294 2071
rect 3478 2068 3497 2071
rect 2142 2058 2161 2061
rect 2174 2058 2201 2061
rect 2314 2058 2321 2061
rect 2426 2058 2433 2061
rect 2542 2061 2545 2068
rect 2526 2058 2545 2061
rect 2958 2058 2974 2061
rect 3226 2058 3233 2061
rect 3454 2058 3470 2061
rect 66 2048 70 2052
rect 110 2048 129 2051
rect 638 2048 646 2051
rect 894 2048 905 2051
rect 1782 2048 1793 2051
rect 1798 2048 1801 2058
rect 1782 2042 1785 2048
rect 98 2038 99 2042
rect 838 2038 862 2041
rect 1746 2038 1747 2042
rect 2677 2038 2678 2042
rect 3506 2038 3507 2042
rect 3710 2038 3718 2041
rect 2434 2028 2435 2032
rect 1234 2018 1235 2022
rect 1258 2018 1259 2022
rect 3402 2018 3403 2022
rect 344 2003 346 2007
rect 350 2003 353 2007
rect 357 2003 360 2007
rect 1360 2003 1362 2007
rect 1366 2003 1369 2007
rect 1373 2003 1376 2007
rect 2384 2003 2386 2007
rect 2390 2003 2393 2007
rect 2397 2003 2400 2007
rect 3408 2003 3410 2007
rect 3414 2003 3417 2007
rect 3421 2003 3424 2007
rect 274 1988 275 1992
rect 594 1988 595 1992
rect 1013 1988 1014 1992
rect 1570 1988 1571 1992
rect 1730 1988 1731 1992
rect 1794 1988 1795 1992
rect 2858 1988 2859 1992
rect 2941 1988 2942 1992
rect 622 1971 625 1981
rect 1634 1978 1635 1982
rect 2330 1978 2331 1982
rect 606 1968 625 1971
rect 1038 1968 1062 1971
rect 1170 1968 1185 1971
rect 1762 1968 1763 1972
rect 3730 1968 3753 1971
rect 66 1958 70 1962
rect 78 1958 97 1961
rect 1054 1958 1065 1961
rect 1054 1952 1058 1954
rect 266 1948 273 1951
rect 554 1948 561 1951
rect 682 1948 689 1951
rect 730 1948 737 1951
rect 1422 1951 1425 1961
rect 1422 1948 1441 1951
rect 1646 1951 1649 1961
rect 2014 1958 2033 1961
rect 2738 1958 2742 1962
rect 3126 1958 3137 1961
rect 1646 1948 1665 1951
rect 1874 1948 1897 1951
rect 1994 1948 2001 1951
rect 2006 1948 2022 1951
rect 2266 1948 2273 1951
rect 2386 1948 2398 1951
rect 2494 1948 2521 1951
rect 2598 1951 2601 1958
rect 2598 1948 2609 1951
rect 2654 1948 2673 1951
rect 2678 1948 2705 1951
rect 3230 1948 3238 1951
rect 3270 1948 3278 1951
rect 3470 1948 3478 1951
rect 310 1941 313 1948
rect 310 1938 321 1941
rect 942 1938 953 1941
rect 1359 1938 1393 1941
rect 1594 1938 1601 1941
rect 2198 1938 2201 1948
rect 2222 1938 2241 1941
rect 2290 1938 2305 1941
rect 2354 1938 2361 1941
rect 2614 1938 2633 1941
rect 3026 1938 3038 1941
rect 3294 1938 3305 1941
rect 3314 1938 3321 1941
rect 3326 1938 3353 1941
rect 3366 1938 3393 1941
rect 3418 1938 3433 1941
rect 3458 1938 3465 1941
rect 3474 1938 3481 1941
rect 3542 1938 3553 1941
rect 3598 1938 3609 1941
rect 2374 1928 2382 1931
rect 2630 1928 2633 1938
rect 3302 1932 3305 1938
rect 3526 1931 3529 1938
rect 3550 1932 3553 1938
rect 3606 1932 3609 1938
rect 3674 1938 3681 1941
rect 3518 1928 3529 1931
rect 3630 1931 3633 1938
rect 3622 1928 3633 1931
rect 1074 1918 1081 1921
rect 1140 1918 1142 1922
rect 1418 1918 1419 1922
rect 3365 1918 3366 1922
rect 3746 1918 3753 1921
rect 848 1903 850 1907
rect 854 1903 857 1907
rect 861 1903 864 1907
rect 1880 1903 1882 1907
rect 1886 1903 1889 1907
rect 1893 1903 1896 1907
rect 2904 1903 2906 1907
rect 2910 1903 2913 1907
rect 2917 1903 2920 1907
rect 666 1888 667 1892
rect 805 1888 806 1892
rect 1229 1888 1230 1892
rect 1594 1888 1595 1892
rect 1618 1888 1619 1892
rect 2370 1888 2371 1892
rect 2946 1888 2947 1892
rect 822 1878 830 1882
rect 2046 1878 2057 1881
rect 822 1872 825 1878
rect 38 1868 57 1871
rect 410 1868 441 1871
rect 1206 1871 1209 1878
rect 1190 1868 1209 1871
rect 2078 1868 2097 1871
rect 2382 1868 2406 1871
rect 2438 1871 2441 1881
rect 3598 1878 3606 1881
rect 2422 1868 2441 1871
rect 2466 1868 2473 1871
rect 2954 1868 2969 1871
rect 3338 1868 3361 1871
rect 3390 1868 3417 1871
rect 3462 1868 3470 1871
rect 3498 1868 3505 1871
rect 2078 1862 2081 1868
rect 246 1852 249 1862
rect 498 1858 505 1861
rect 750 1858 769 1861
rect 1038 1858 1062 1861
rect 1094 1858 1102 1861
rect 1110 1858 1137 1861
rect 1166 1858 1185 1861
rect 1262 1858 1289 1861
rect 1298 1858 1313 1861
rect 1502 1858 1510 1861
rect 1910 1858 1929 1861
rect 1942 1858 1969 1861
rect 1974 1858 2001 1861
rect 2462 1858 2470 1861
rect 2546 1858 2561 1861
rect 2766 1858 2790 1861
rect 2846 1861 2849 1868
rect 2846 1858 2857 1861
rect 2862 1858 2870 1861
rect 3186 1858 3193 1861
rect 3238 1858 3246 1861
rect 3414 1861 3417 1868
rect 3638 1862 3641 1871
rect 3414 1858 3433 1861
rect 518 1848 526 1851
rect 766 1848 769 1858
rect 1478 1852 1482 1854
rect 958 1848 966 1851
rect 1150 1848 1169 1851
rect 1258 1848 1262 1852
rect 1558 1848 1569 1851
rect 1926 1848 1929 1858
rect 2794 1848 2798 1852
rect 2934 1851 2937 1858
rect 2926 1848 2937 1851
rect 2954 1848 2961 1851
rect 3170 1848 3174 1852
rect 1558 1842 1562 1844
rect 658 1838 665 1841
rect 3654 1838 3662 1841
rect 566 1828 569 1838
rect 781 1818 782 1822
rect 2501 1818 2502 1822
rect 2562 1818 2563 1822
rect 3514 1818 3515 1822
rect 344 1803 346 1807
rect 350 1803 353 1807
rect 357 1803 360 1807
rect 1360 1803 1362 1807
rect 1366 1803 1369 1807
rect 1373 1803 1376 1807
rect 2384 1803 2386 1807
rect 2390 1803 2393 1807
rect 2397 1803 2400 1807
rect 3408 1803 3410 1807
rect 3414 1803 3417 1807
rect 3421 1803 3424 1807
rect 458 1788 459 1792
rect 874 1788 889 1791
rect 1597 1788 1598 1792
rect 294 1768 305 1771
rect 982 1768 990 1771
rect 1565 1768 1566 1772
rect 1930 1768 1931 1772
rect 2266 1768 2273 1771
rect 2693 1768 2694 1772
rect 2882 1768 2883 1772
rect 3622 1771 3625 1781
rect 3622 1768 3657 1771
rect 302 1758 305 1768
rect 1010 1758 1014 1762
rect 1626 1758 1630 1762
rect 1942 1758 1953 1761
rect 2466 1758 2470 1762
rect 22 1748 41 1751
rect 362 1748 377 1751
rect 474 1748 481 1751
rect 542 1748 550 1751
rect 658 1748 665 1751
rect 782 1748 790 1751
rect 1002 1748 1009 1751
rect 1566 1748 1574 1751
rect 1618 1748 1625 1751
rect 2030 1748 2041 1751
rect 2138 1748 2153 1751
rect 2586 1748 2593 1751
rect 2642 1748 2649 1751
rect 2758 1748 2785 1751
rect 2798 1751 2801 1761
rect 2894 1758 2921 1761
rect 2798 1748 2817 1751
rect 2978 1748 2985 1751
rect 3038 1751 3042 1752
rect 3022 1748 3042 1751
rect 3158 1751 3162 1754
rect 3142 1748 3162 1751
rect 3246 1748 3265 1751
rect 3318 1748 3329 1751
rect 3358 1748 3377 1751
rect 3726 1751 3730 1754
rect 3726 1748 3745 1751
rect 334 1738 345 1741
rect 862 1738 886 1741
rect 950 1741 953 1748
rect 950 1738 961 1741
rect 1054 1738 1062 1741
rect 1458 1738 1465 1741
rect 1990 1738 2006 1741
rect 2034 1738 2049 1741
rect 2066 1738 2073 1741
rect 2486 1738 2489 1748
rect 2938 1738 2961 1741
rect 3494 1738 3513 1741
rect 3582 1738 3593 1741
rect 334 1732 337 1738
rect 3590 1732 3593 1738
rect 390 1728 401 1731
rect 2134 1728 2142 1731
rect 2214 1728 2233 1731
rect 1253 1718 1254 1722
rect 1474 1718 1475 1722
rect 1901 1718 1902 1722
rect 3406 1718 3422 1721
rect 3674 1718 3676 1722
rect 3710 1718 3718 1721
rect 3754 1718 3756 1722
rect 848 1703 850 1707
rect 854 1703 857 1707
rect 861 1703 864 1707
rect 1880 1703 1882 1707
rect 1886 1703 1889 1707
rect 1893 1703 1896 1707
rect 2904 1703 2906 1707
rect 2910 1703 2913 1707
rect 2917 1703 2920 1707
rect 581 1688 582 1692
rect 1210 1688 1217 1691
rect 1541 1688 1542 1692
rect 3082 1688 3083 1692
rect 3125 1688 3126 1692
rect 3253 1688 3254 1692
rect 3746 1688 3748 1692
rect 370 1678 385 1681
rect 1718 1678 1729 1681
rect 1798 1678 1817 1681
rect 1950 1678 1969 1681
rect 2066 1678 2073 1681
rect 2342 1678 2358 1681
rect 2742 1678 2753 1681
rect 2934 1678 2945 1681
rect 3290 1678 3297 1681
rect 3434 1678 3441 1681
rect 3558 1678 3569 1681
rect 3638 1678 3649 1681
rect 690 1668 697 1671
rect 302 1658 305 1668
rect 370 1658 377 1661
rect 790 1661 793 1671
rect 1422 1668 1433 1671
rect 1518 1671 1521 1678
rect 1726 1672 1729 1678
rect 1510 1668 1521 1671
rect 1738 1668 1745 1671
rect 1822 1671 1825 1678
rect 3566 1672 3569 1678
rect 3646 1672 3649 1678
rect 1822 1668 1833 1671
rect 1878 1668 1902 1671
rect 2602 1668 2609 1671
rect 2842 1668 2857 1671
rect 2874 1668 2881 1671
rect 2982 1668 3001 1671
rect 3062 1668 3070 1671
rect 3090 1668 3105 1671
rect 3406 1668 3438 1671
rect 3446 1668 3465 1671
rect 3502 1668 3521 1671
rect 778 1658 793 1661
rect 958 1658 966 1661
rect 998 1658 1017 1661
rect 1206 1658 1209 1668
rect 1278 1658 1297 1661
rect 1386 1658 1409 1661
rect 1446 1658 1473 1661
rect 1719 1658 1737 1661
rect 1878 1661 1881 1668
rect 2982 1662 2985 1668
rect 1874 1658 1881 1661
rect 2082 1658 2089 1661
rect 2806 1658 2814 1661
rect 2862 1658 2870 1661
rect 3510 1658 3518 1661
rect 3602 1658 3609 1661
rect 3658 1658 3665 1661
rect 574 1648 577 1658
rect 814 1648 822 1651
rect 1014 1648 1017 1658
rect 1142 1652 1146 1654
rect 1294 1648 1297 1658
rect 1302 1648 1321 1651
rect 1526 1648 1537 1651
rect 1870 1648 1886 1651
rect 2022 1648 2033 1651
rect 2598 1648 2609 1651
rect 678 1642 682 1644
rect 622 1638 641 1641
rect 1094 1641 1098 1644
rect 1086 1638 1098 1641
rect 1858 1638 1859 1642
rect 638 1628 641 1638
rect 2701 1618 2702 1622
rect 344 1603 346 1607
rect 350 1603 353 1607
rect 357 1603 360 1607
rect 1360 1603 1362 1607
rect 1366 1603 1369 1607
rect 1373 1603 1376 1607
rect 2384 1603 2386 1607
rect 2390 1603 2393 1607
rect 2397 1603 2400 1607
rect 3408 1603 3410 1607
rect 3414 1603 3417 1607
rect 3421 1603 3424 1607
rect 970 1588 971 1592
rect 1493 1588 1494 1592
rect 3538 1588 3539 1592
rect 474 1578 475 1582
rect 1166 1568 1177 1571
rect 2898 1568 2899 1572
rect 3622 1568 3633 1571
rect 1166 1562 1169 1568
rect 3622 1562 3625 1568
rect 742 1558 750 1561
rect 454 1548 473 1551
rect 522 1548 537 1551
rect 722 1548 729 1551
rect 734 1548 742 1551
rect 774 1548 785 1551
rect 962 1548 969 1551
rect 1478 1551 1481 1561
rect 3010 1558 3014 1562
rect 3554 1558 3561 1561
rect 1462 1548 1481 1551
rect 1846 1548 1857 1551
rect 1890 1548 1905 1551
rect 590 1538 593 1548
rect 1982 1542 1985 1551
rect 2574 1548 2593 1551
rect 2598 1548 2614 1551
rect 2882 1548 2897 1551
rect 3014 1548 3022 1551
rect 3038 1548 3046 1551
rect 3062 1548 3078 1551
rect 2318 1538 2326 1541
rect 2534 1538 2553 1541
rect 3022 1538 3041 1541
rect 3478 1538 3486 1541
rect 3518 1538 3526 1541
rect 1806 1528 1825 1531
rect 2294 1528 2297 1538
rect 2550 1528 2553 1538
rect 3102 1528 3113 1531
rect 3546 1528 3553 1531
rect 3558 1528 3569 1531
rect 3642 1528 3649 1531
rect 309 1518 310 1522
rect 1093 1518 1094 1522
rect 1117 1518 1118 1522
rect 1141 1518 1142 1522
rect 3309 1518 3310 1522
rect 3421 1518 3422 1522
rect 848 1503 850 1507
rect 854 1503 857 1507
rect 861 1503 864 1507
rect 1880 1503 1882 1507
rect 1886 1503 1889 1507
rect 1893 1503 1896 1507
rect 2904 1503 2906 1507
rect 2910 1503 2913 1507
rect 2917 1503 2920 1507
rect 1026 1488 1027 1492
rect 1882 1488 1897 1491
rect 342 1478 366 1481
rect 1838 1478 1849 1481
rect 2534 1478 2545 1481
rect 3058 1478 3065 1481
rect 3118 1478 3129 1481
rect 3246 1478 3257 1481
rect 3286 1478 3294 1481
rect 3562 1478 3569 1481
rect 3654 1478 3662 1481
rect 3118 1472 3121 1478
rect 3246 1472 3249 1478
rect 814 1462 817 1471
rect 874 1468 897 1471
rect 1110 1468 1134 1471
rect 1154 1468 1161 1471
rect 1198 1468 1209 1471
rect 1334 1468 1350 1471
rect 414 1458 433 1461
rect 526 1458 534 1461
rect 910 1458 918 1461
rect 970 1458 985 1461
rect 1030 1461 1033 1468
rect 1198 1462 1201 1468
rect 1030 1458 1041 1461
rect 1078 1458 1086 1461
rect 1766 1458 1785 1461
rect 2350 1461 2353 1468
rect 2322 1458 2329 1461
rect 2342 1458 2353 1461
rect 2382 1458 2425 1461
rect 2430 1458 2457 1461
rect 2614 1461 2617 1468
rect 2998 1468 3006 1471
rect 3062 1468 3073 1471
rect 3102 1468 3110 1471
rect 3150 1468 3161 1471
rect 3382 1468 3390 1471
rect 3498 1468 3521 1471
rect 3574 1468 3593 1471
rect 3630 1468 3638 1471
rect 3062 1462 3065 1468
rect 3158 1462 3161 1468
rect 2614 1458 2625 1461
rect 2670 1458 2678 1461
rect 2702 1458 2729 1461
rect 2830 1458 2846 1461
rect 2902 1458 2926 1461
rect 3018 1458 3025 1461
rect 3238 1458 3249 1461
rect 3594 1458 3601 1461
rect 18 1448 25 1451
rect 402 1448 407 1452
rect 846 1448 849 1458
rect 1074 1448 1078 1452
rect 1782 1448 1785 1458
rect 2342 1448 2345 1458
rect 2402 1448 2417 1451
rect 2858 1448 2862 1452
rect 3470 1448 3481 1451
rect 726 1442 730 1444
rect 1030 1442 1034 1444
rect 2669 1438 2670 1442
rect 2797 1438 2798 1442
rect 2701 1418 2702 1422
rect 2762 1418 2763 1422
rect 2970 1418 2971 1422
rect 3458 1418 3459 1422
rect 344 1403 346 1407
rect 350 1403 353 1407
rect 357 1403 360 1407
rect 1360 1403 1362 1407
rect 1366 1403 1369 1407
rect 1373 1403 1376 1407
rect 2384 1403 2386 1407
rect 2390 1403 2393 1407
rect 2397 1403 2400 1407
rect 3408 1403 3410 1407
rect 3414 1403 3417 1407
rect 3421 1403 3424 1407
rect 258 1388 259 1392
rect 522 1388 523 1392
rect 1565 1388 1566 1392
rect 1714 1388 1715 1392
rect 1789 1388 1790 1392
rect 1821 1388 1822 1392
rect 3546 1388 3547 1392
rect 478 1368 486 1371
rect 578 1368 579 1372
rect 710 1371 713 1381
rect 3702 1372 3705 1381
rect 694 1368 713 1371
rect 1650 1368 1651 1372
rect 2117 1368 2118 1372
rect 2853 1368 2854 1372
rect 790 1358 801 1361
rect 62 1348 81 1351
rect 250 1348 257 1351
rect 494 1348 513 1351
rect 834 1348 841 1351
rect 910 1348 918 1351
rect 990 1348 998 1351
rect 1414 1351 1417 1361
rect 1398 1348 1417 1351
rect 1442 1348 1457 1351
rect 1598 1351 1601 1361
rect 1570 1348 1585 1351
rect 1598 1348 1617 1351
rect 1662 1351 1665 1361
rect 1662 1348 1681 1351
rect 1822 1348 1849 1351
rect 2102 1351 2105 1361
rect 2086 1348 2105 1351
rect 2118 1348 2145 1351
rect 2150 1348 2177 1351
rect 2270 1351 2273 1361
rect 2270 1348 2281 1351
rect 2310 1348 2337 1351
rect 2342 1348 2369 1351
rect 2438 1351 2441 1361
rect 2906 1358 2921 1361
rect 3446 1358 3454 1361
rect 2402 1348 2417 1351
rect 2422 1348 2441 1351
rect 2454 1348 2481 1351
rect 2486 1348 2513 1351
rect 2810 1348 2817 1351
rect 2822 1348 2838 1351
rect 3094 1348 3102 1351
rect 510 1342 513 1348
rect 542 1338 556 1341
rect 590 1338 593 1348
rect 1410 1338 1417 1341
rect 1470 1338 1481 1341
rect 1582 1338 1585 1348
rect 1734 1338 1742 1341
rect 2198 1341 2201 1348
rect 2278 1342 2281 1348
rect 2198 1338 2209 1341
rect 2946 1338 2961 1341
rect 3062 1341 3065 1348
rect 3230 1342 3233 1351
rect 3294 1348 3313 1351
rect 3602 1348 3609 1351
rect 3062 1338 3081 1341
rect 3154 1338 3161 1341
rect 3246 1338 3273 1341
rect 3286 1338 3294 1341
rect 542 1332 545 1338
rect 1366 1328 1374 1331
rect 1526 1331 1529 1338
rect 3614 1332 3617 1351
rect 3650 1348 3657 1351
rect 3766 1348 3774 1351
rect 3670 1338 3678 1341
rect 1526 1328 1537 1331
rect 1878 1328 1902 1331
rect 2894 1328 2921 1331
rect 854 1318 870 1321
rect 938 1318 939 1322
rect 3138 1318 3139 1322
rect 848 1303 850 1307
rect 854 1303 857 1307
rect 861 1303 864 1307
rect 1880 1303 1882 1307
rect 1886 1303 1889 1307
rect 1893 1303 1896 1307
rect 2904 1303 2906 1307
rect 2910 1303 2913 1307
rect 2917 1303 2920 1307
rect 3578 1288 3579 1292
rect 1422 1278 1441 1281
rect 190 1268 201 1271
rect 206 1268 225 1271
rect 1078 1268 1097 1271
rect 1390 1271 1393 1278
rect 1390 1268 1401 1271
rect 1486 1268 1505 1271
rect 1618 1268 1625 1271
rect 2022 1271 2025 1281
rect 2262 1278 2273 1281
rect 3742 1278 3750 1282
rect 3742 1272 3745 1278
rect 2022 1268 2041 1271
rect 2378 1268 2401 1271
rect 2486 1268 2505 1271
rect 2590 1268 2609 1271
rect 2914 1268 2921 1271
rect 3118 1268 3126 1271
rect 3130 1268 3137 1271
rect 3390 1268 3398 1271
rect 3694 1268 3721 1271
rect 222 1262 226 1264
rect 2486 1262 2489 1268
rect 510 1258 529 1261
rect 1046 1258 1065 1261
rect 1110 1258 1118 1261
rect 1462 1258 1473 1261
rect 1494 1258 1502 1261
rect 2014 1258 2022 1261
rect 2374 1258 2382 1261
rect 2426 1258 2433 1261
rect 2886 1258 2902 1261
rect 2962 1258 2969 1261
rect 2978 1258 2993 1261
rect 3150 1258 3177 1261
rect 3194 1258 3201 1261
rect 3242 1258 3250 1261
rect 3358 1258 3369 1261
rect 3398 1258 3417 1261
rect 3518 1258 3537 1261
rect 510 1248 513 1258
rect 538 1248 545 1251
rect 1062 1248 1065 1258
rect 1574 1248 1585 1251
rect 2630 1248 2638 1251
rect 2842 1238 2843 1242
rect 2618 1228 2619 1232
rect 994 1218 995 1222
rect 2317 1218 2318 1222
rect 2994 1218 2995 1222
rect 3069 1218 3070 1222
rect 3178 1218 3179 1222
rect 344 1203 346 1207
rect 350 1203 353 1207
rect 357 1203 360 1207
rect 1360 1203 1362 1207
rect 1366 1203 1369 1207
rect 1373 1203 1376 1207
rect 2384 1203 2386 1207
rect 2390 1203 2393 1207
rect 2397 1203 2400 1207
rect 3408 1203 3410 1207
rect 3414 1203 3417 1207
rect 3421 1203 3424 1207
rect 221 1188 222 1192
rect 250 1188 251 1192
rect 1058 1188 1059 1192
rect 2301 1188 2302 1192
rect 3106 1188 3107 1192
rect 3221 1188 3222 1192
rect 838 1171 841 1181
rect 1917 1178 1918 1182
rect 3554 1178 3555 1182
rect 822 1168 841 1171
rect 3730 1168 3731 1172
rect 910 1166 914 1168
rect 18 1158 25 1161
rect 167 1148 174 1151
rect 206 1151 209 1161
rect 1018 1158 1025 1161
rect 198 1148 209 1151
rect 254 1148 262 1151
rect 398 1148 422 1151
rect 790 1148 806 1151
rect 874 1148 889 1151
rect 910 1148 921 1151
rect 1366 1151 1369 1161
rect 1570 1158 1574 1162
rect 1582 1158 1593 1161
rect 1366 1148 1401 1151
rect 1526 1148 1534 1151
rect 1638 1148 1646 1151
rect 1862 1151 1865 1158
rect 1862 1148 1873 1151
rect 2390 1148 2414 1151
rect 2558 1148 2569 1151
rect 2846 1151 2849 1161
rect 3506 1158 3513 1161
rect 2830 1148 2849 1151
rect 2906 1148 2929 1151
rect 2934 1148 2961 1151
rect 910 1142 913 1148
rect 3006 1142 3009 1151
rect 3270 1148 3281 1151
rect 3310 1148 3329 1151
rect 3546 1148 3553 1151
rect 3570 1148 3585 1151
rect 230 1138 241 1141
rect 238 1132 241 1138
rect 254 1138 265 1141
rect 350 1138 358 1141
rect 362 1138 377 1141
rect 562 1138 569 1141
rect 1134 1138 1145 1141
rect 1498 1138 1513 1141
rect 1642 1138 1649 1141
rect 2402 1138 2433 1141
rect 2590 1138 2609 1141
rect 2974 1138 2982 1141
rect 2990 1138 3006 1141
rect 3438 1138 3449 1141
rect 3478 1138 3481 1148
rect 3650 1138 3665 1141
rect 3714 1138 3721 1141
rect 254 1132 257 1138
rect 166 1128 185 1131
rect 1150 1128 1158 1131
rect 1486 1128 1505 1131
rect 1630 1128 1638 1131
rect 1862 1128 1865 1138
rect 2342 1128 2353 1131
rect 2590 1128 2593 1138
rect 3446 1132 3449 1138
rect 2630 1128 2638 1131
rect 3078 1128 3086 1131
rect 3150 1128 3158 1131
rect 3174 1128 3185 1131
rect 3398 1128 3414 1131
rect 485 1118 486 1122
rect 1010 1118 1011 1122
rect 1029 1118 1030 1122
rect 1366 1118 1382 1121
rect 1429 1118 1430 1122
rect 2885 1118 2886 1122
rect 848 1103 850 1107
rect 854 1103 857 1107
rect 861 1103 864 1107
rect 1880 1103 1882 1107
rect 1886 1103 1889 1107
rect 1893 1103 1896 1107
rect 2904 1103 2906 1107
rect 2910 1103 2913 1107
rect 2917 1103 2920 1107
rect 1634 1088 1635 1092
rect 1514 1078 1521 1081
rect 250 1068 257 1071
rect 958 1062 961 1071
rect 1406 1068 1417 1071
rect 1474 1068 1481 1071
rect 1566 1071 1569 1081
rect 1550 1068 1569 1071
rect 1614 1068 1622 1071
rect 1638 1068 1649 1071
rect 1766 1071 1769 1081
rect 1750 1068 1769 1071
rect 1975 1068 1993 1071
rect 2090 1068 2113 1071
rect 2174 1071 2177 1078
rect 2174 1068 2185 1071
rect 2214 1068 2222 1071
rect 2294 1071 2297 1081
rect 3058 1078 3065 1081
rect 2278 1068 2297 1071
rect 2798 1068 2806 1071
rect 2866 1068 2881 1071
rect 3134 1068 3142 1071
rect 3366 1068 3385 1071
rect 3494 1068 3505 1071
rect 3518 1068 3545 1071
rect 1638 1062 1641 1068
rect 3502 1062 3505 1068
rect 318 1058 326 1061
rect 718 1058 726 1061
rect 1350 1058 1374 1061
rect 1430 1058 1449 1061
rect 1790 1058 1798 1061
rect 2318 1058 2329 1061
rect 2362 1058 2369 1061
rect 2618 1058 2625 1061
rect 2834 1058 2857 1061
rect 2894 1058 2918 1061
rect 3002 1058 3009 1061
rect 3186 1058 3193 1061
rect 3350 1058 3358 1061
rect 3374 1058 3382 1061
rect 3606 1058 3622 1061
rect 246 1048 254 1051
rect 310 1042 313 1051
rect 330 1048 361 1051
rect 726 1048 745 1051
rect 1722 1048 1726 1052
rect 2018 1048 2022 1052
rect 2370 1048 2374 1052
rect 2382 1048 2409 1051
rect 2610 1048 2617 1051
rect 2722 1048 2726 1052
rect 2734 1048 2737 1058
rect 3074 1048 3081 1051
rect 2933 1028 2934 1032
rect 3634 1028 3635 1032
rect 1133 1018 1134 1022
rect 1253 1018 1254 1022
rect 1690 1018 1691 1022
rect 2053 1018 2054 1022
rect 2514 1018 2515 1022
rect 2690 1018 2691 1022
rect 3050 1018 3051 1022
rect 3205 1018 3206 1022
rect 3394 1018 3395 1022
rect 344 1003 346 1007
rect 350 1003 353 1007
rect 357 1003 360 1007
rect 1360 1003 1362 1007
rect 1366 1003 1369 1007
rect 1373 1003 1376 1007
rect 2384 1003 2386 1007
rect 2390 1003 2393 1007
rect 2397 1003 2400 1007
rect 3408 1003 3410 1007
rect 3414 1003 3417 1007
rect 3421 1003 3424 1007
rect 1578 988 1579 992
rect 2938 988 2939 992
rect 242 978 243 982
rect 3494 972 3497 981
rect 3582 972 3585 981
rect 2674 968 2681 971
rect 50 958 57 961
rect 254 958 262 961
rect 278 958 286 961
rect 222 948 241 951
rect 346 948 361 951
rect 414 951 417 961
rect 930 958 937 961
rect 398 948 417 951
rect 502 948 513 951
rect 922 948 945 951
rect 1646 948 1654 951
rect 1702 951 1705 961
rect 1702 948 1721 951
rect 1918 948 1937 951
rect 2318 948 2345 951
rect 2350 948 2377 951
rect 2594 948 2601 951
rect 2750 948 2769 951
rect 474 938 481 941
rect 558 938 566 941
rect 1166 938 1193 941
rect 1198 938 1217 941
rect 1626 938 1633 941
rect 1758 938 1766 941
rect 1898 938 1905 941
rect 2278 938 2281 948
rect 2450 938 2457 941
rect 2750 938 2753 948
rect 2814 938 2817 958
rect 2894 948 2918 951
rect 3022 951 3026 954
rect 3006 948 3026 951
rect 3346 948 3353 951
rect 3414 948 3457 951
rect 3690 948 3697 951
rect 3742 948 3761 951
rect 3222 938 3238 941
rect 3298 938 3305 941
rect 3366 938 3369 948
rect 3710 938 3721 941
rect 2222 932 2225 938
rect 570 928 577 931
rect 2218 928 2225 932
rect 2850 928 2854 932
rect 3286 931 3289 938
rect 3278 928 3289 931
rect 274 918 275 922
rect 549 918 550 922
rect 1674 918 1675 922
rect 2661 918 2662 922
rect 3642 918 3643 922
rect 848 903 850 907
rect 854 903 857 907
rect 861 903 864 907
rect 1880 903 1882 907
rect 1886 903 1889 907
rect 1893 903 1896 907
rect 2904 903 2906 907
rect 2910 903 2913 907
rect 2917 903 2920 907
rect 1861 888 1862 892
rect 1922 888 1923 892
rect 2378 888 2379 892
rect 2402 888 2409 891
rect 1314 878 1337 881
rect 1614 878 1633 881
rect 1694 878 1705 881
rect 2574 878 2593 881
rect 2762 878 2769 882
rect 3414 878 3441 881
rect 3534 878 3545 881
rect 590 876 594 878
rect 482 868 489 871
rect 514 868 529 871
rect 1270 868 1278 871
rect 1534 862 1537 871
rect 1670 868 1689 871
rect 1710 868 1721 871
rect 1746 868 1761 871
rect 1906 868 1921 871
rect 1934 868 1950 871
rect 2486 871 2489 878
rect 2766 872 2769 878
rect 2486 868 2505 871
rect 2594 868 2601 871
rect 2946 868 2953 871
rect 3198 868 3206 871
rect 3238 868 3246 871
rect 3262 868 3270 871
rect 3310 868 3318 871
rect 3390 868 3398 871
rect 3562 868 3569 871
rect 3654 868 3665 871
rect 3730 868 3737 871
rect 1710 862 1713 868
rect 3662 862 3665 868
rect 190 858 209 861
rect 478 858 486 861
rect 506 858 521 861
rect 1554 858 1577 861
rect 2318 858 2337 861
rect 2486 858 2494 861
rect 2690 858 2697 861
rect 2942 858 2950 861
rect 3242 858 3249 861
rect 3622 858 3630 861
rect 18 848 25 851
rect 486 848 489 858
rect 1246 848 1257 851
rect 1514 848 1518 852
rect 1786 848 1790 852
rect 1890 848 1897 851
rect 2334 848 2337 858
rect 2394 848 2409 851
rect 2714 848 2721 851
rect 2870 848 2881 851
rect 3114 848 3118 852
rect 3178 838 3179 842
rect 1661 828 1662 832
rect 3085 828 3086 832
rect 474 818 475 822
rect 562 818 563 822
rect 1117 818 1118 822
rect 2482 818 2483 822
rect 2530 818 2531 822
rect 2554 818 2555 822
rect 2698 818 2699 822
rect 2733 818 2734 822
rect 2826 818 2827 822
rect 2858 818 2859 822
rect 3146 818 3147 822
rect 3229 818 3230 822
rect 344 803 346 807
rect 350 803 353 807
rect 357 803 360 807
rect 1360 803 1362 807
rect 1366 803 1369 807
rect 1373 803 1376 807
rect 2384 803 2386 807
rect 2390 803 2393 807
rect 2397 803 2400 807
rect 3408 803 3410 807
rect 3414 803 3417 807
rect 3421 803 3424 807
rect 282 788 283 792
rect 394 788 395 792
rect 794 788 795 792
rect 2346 788 2347 792
rect 3434 788 3435 792
rect 3522 788 3523 792
rect 3586 788 3587 792
rect 189 778 190 782
rect 310 768 318 771
rect 365 768 366 772
rect 822 771 825 781
rect 1690 778 1691 782
rect 806 768 825 771
rect 3730 768 3731 772
rect 34 748 41 751
rect 102 748 113 751
rect 1222 751 1225 758
rect 1198 748 1217 751
rect 1222 748 1233 751
rect 1522 748 1529 751
rect 1570 748 1585 751
rect 1622 748 1630 751
rect 2086 751 2089 761
rect 2766 758 2777 761
rect 2978 758 2982 762
rect 2990 758 3001 761
rect 2070 748 2089 751
rect 2266 748 2273 751
rect 2458 748 2465 751
rect 2470 748 2486 751
rect 2758 748 2766 751
rect 3062 748 3073 751
rect 3146 748 3153 751
rect 126 738 134 741
rect 146 738 153 741
rect 242 738 249 741
rect 318 738 329 741
rect 502 741 505 748
rect 502 738 521 741
rect 1246 738 1265 741
rect 1270 738 1289 741
rect 1514 738 1521 741
rect 1590 738 1606 741
rect 1662 738 1681 741
rect 1758 738 1774 741
rect 1806 741 1809 748
rect 1806 738 1817 741
rect 2082 738 2089 741
rect 2154 738 2161 741
rect 2286 738 2294 741
rect 2790 738 2798 741
rect 3198 741 3201 751
rect 3330 748 3337 751
rect 3366 748 3382 751
rect 3414 748 3433 751
rect 3470 748 3478 751
rect 3646 748 3657 751
rect 3722 748 3729 751
rect 3138 738 3145 741
rect 3182 738 3201 741
rect 3294 738 3302 741
rect 3414 741 3417 748
rect 3654 742 3657 748
rect 3390 738 3417 741
rect 3670 738 3678 741
rect 1270 732 1273 738
rect 374 728 382 731
rect 466 728 470 732
rect 530 728 545 731
rect 1646 728 1657 731
rect 2950 728 2958 731
rect 2898 718 2913 721
rect 3754 718 3756 722
rect 848 703 850 707
rect 854 703 857 707
rect 861 703 864 707
rect 1880 703 1882 707
rect 1886 703 1889 707
rect 1893 703 1896 707
rect 2904 703 2906 707
rect 2910 703 2913 707
rect 2917 703 2920 707
rect 554 688 556 692
rect 2485 688 2486 692
rect 2802 688 2803 692
rect 2842 688 2843 692
rect 2901 688 2902 692
rect 2986 688 2987 692
rect 3069 688 3070 692
rect 3466 688 3467 692
rect 3709 688 3710 692
rect 198 678 206 681
rect 494 678 505 681
rect 1318 678 1326 682
rect 1374 678 1398 681
rect 1470 678 1478 681
rect 1550 678 1561 681
rect 2714 678 2721 681
rect 2954 678 2961 681
rect 3758 678 3766 682
rect 190 668 198 671
rect 398 671 401 678
rect 1318 672 1321 678
rect 3758 672 3761 678
rect 342 668 369 671
rect 398 668 409 671
rect 202 658 209 661
rect 214 658 233 661
rect 534 661 537 671
rect 830 668 865 671
rect 1270 668 1297 671
rect 1342 668 1350 671
rect 1378 668 1409 671
rect 1526 668 1545 671
rect 1566 668 1577 671
rect 1622 668 1630 671
rect 1634 668 1641 671
rect 1823 668 1841 671
rect 1858 668 1865 671
rect 522 658 537 661
rect 1014 658 1017 668
rect 1566 662 1569 668
rect 2022 662 2025 671
rect 2110 668 2129 671
rect 2382 668 2398 671
rect 2518 668 2526 671
rect 2754 668 2761 671
rect 2774 668 2782 671
rect 2850 668 2865 671
rect 3622 668 3630 671
rect 1846 658 1865 661
rect 1878 658 1921 661
rect 1990 658 1998 661
rect 2070 658 2097 661
rect 2126 658 2134 661
rect 2374 658 2417 661
rect 2422 658 2430 661
rect 3054 658 3062 661
rect 3082 658 3089 661
rect 3294 661 3297 668
rect 3294 658 3305 661
rect 3434 658 3441 661
rect 3670 658 3689 661
rect 3718 658 3729 661
rect 18 648 25 651
rect 230 648 233 658
rect 1638 651 1641 658
rect 1638 648 1649 651
rect 1862 648 1865 658
rect 1898 648 1913 651
rect 2806 648 2817 651
rect 3282 648 3286 652
rect 2814 638 2822 641
rect 2974 641 2977 648
rect 2966 638 2977 641
rect 450 618 451 622
rect 1461 618 1462 622
rect 1490 618 1491 622
rect 2946 618 2947 622
rect 3205 618 3206 622
rect 344 603 346 607
rect 350 603 353 607
rect 357 603 360 607
rect 1360 603 1362 607
rect 1366 603 1369 607
rect 1373 603 1376 607
rect 2384 603 2386 607
rect 2390 603 2393 607
rect 2397 603 2400 607
rect 3408 603 3410 607
rect 3414 603 3417 607
rect 3421 603 3424 607
rect 3682 588 3683 592
rect 3754 588 3755 592
rect 3173 578 3174 582
rect 18 558 25 561
rect 262 548 278 551
rect 294 548 302 551
rect 426 548 449 551
rect 530 548 542 551
rect 1214 551 1217 558
rect 1190 548 1209 551
rect 1214 548 1225 551
rect 1526 548 1534 551
rect 302 538 321 541
rect 326 538 358 541
rect 426 538 441 541
rect 814 538 822 541
rect 1062 538 1089 541
rect 1130 538 1137 541
rect 1238 538 1257 541
rect 1406 538 1425 541
rect 1510 541 1513 548
rect 1622 542 1625 551
rect 1706 548 1713 551
rect 1918 551 1921 561
rect 2222 558 2230 561
rect 2706 558 2710 562
rect 1902 548 1921 551
rect 1934 548 1961 551
rect 1966 548 1993 551
rect 2094 548 2102 551
rect 2254 548 2262 551
rect 2442 548 2465 551
rect 2854 548 2862 551
rect 2958 548 2966 551
rect 2998 548 3006 551
rect 3206 548 3214 551
rect 3374 551 3377 561
rect 3374 548 3393 551
rect 3478 548 3486 551
rect 3558 548 3566 551
rect 3746 548 3753 551
rect 1502 538 1513 541
rect 1518 538 1537 541
rect 1638 538 1646 541
rect 1678 538 1686 541
rect 1890 538 1897 541
rect 1914 538 1921 541
rect 2066 538 2081 541
rect 2102 538 2105 548
rect 2510 538 2518 541
rect 2826 538 2841 541
rect 2978 538 2985 541
rect 3058 538 3065 541
rect 3098 538 3105 541
rect 3598 538 3601 548
rect 3718 541 3721 548
rect 3702 538 3721 541
rect 326 528 329 538
rect 482 528 489 531
rect 2934 528 2945 531
rect 3246 528 3257 531
rect 3310 528 3321 531
rect 3446 531 3449 538
rect 3438 528 3449 531
rect 3510 531 3513 538
rect 3502 528 3513 531
rect 1021 518 1022 522
rect 1122 518 1123 522
rect 1357 518 1358 522
rect 1602 518 1603 522
rect 2058 518 2059 522
rect 2818 518 2819 522
rect 848 503 850 507
rect 854 503 857 507
rect 861 503 864 507
rect 1880 503 1882 507
rect 1886 503 1889 507
rect 1893 503 1896 507
rect 2904 503 2906 507
rect 2910 503 2913 507
rect 2917 503 2920 507
rect 202 488 204 492
rect 405 488 406 492
rect 1106 488 1107 492
rect 2613 488 2614 492
rect 438 478 449 481
rect 462 478 473 481
rect 866 478 873 481
rect 1178 478 1179 482
rect 3678 478 3689 481
rect 3750 478 3766 481
rect 446 472 449 478
rect 262 468 273 471
rect 326 468 337 471
rect 414 468 433 471
rect 462 468 473 471
rect 326 462 329 468
rect 414 462 417 468
rect 462 462 465 468
rect 822 462 825 471
rect 878 468 889 471
rect 1202 468 1217 471
rect 1302 468 1321 471
rect 1386 468 1401 471
rect 1822 468 1830 471
rect 1982 471 1985 478
rect 1974 468 1985 471
rect 2314 468 2321 471
rect 2466 468 2473 471
rect 2774 468 2782 471
rect 298 458 313 461
rect 442 458 449 461
rect 522 458 529 461
rect 838 458 881 461
rect 1210 458 1217 461
rect 1318 461 1321 468
rect 1314 458 1321 461
rect 1430 458 1433 468
rect 1494 458 1513 461
rect 1750 458 1769 461
rect 1902 458 1929 461
rect 1934 458 1961 461
rect 2238 458 2265 461
rect 2418 458 2425 461
rect 2430 458 2438 461
rect 2658 458 2673 461
rect 2806 458 2814 461
rect 2842 458 2849 461
rect 2886 458 2921 461
rect 3006 458 3025 461
rect 3226 458 3233 461
rect 3246 461 3249 471
rect 3598 471 3601 478
rect 3590 468 3601 471
rect 3686 468 3697 471
rect 3686 462 3689 468
rect 3246 458 3265 461
rect 3286 458 3313 461
rect 3326 458 3345 461
rect 3706 458 3713 461
rect 1494 456 1498 458
rect 1750 452 1753 458
rect 2182 448 2193 451
rect 2706 448 2710 452
rect 2802 448 2806 452
rect 2918 448 2921 458
rect 2962 448 2966 452
rect 3006 448 3009 458
rect 3326 448 3329 458
rect 1110 442 1114 444
rect 530 438 531 442
rect 806 438 826 441
rect 1358 438 1382 441
rect 1502 441 1506 444
rect 1490 438 1506 441
rect 806 428 809 438
rect 2645 428 2646 432
rect 498 418 499 422
rect 562 418 563 422
rect 2170 418 2171 422
rect 2237 418 2238 422
rect 2365 418 2366 422
rect 2674 418 2675 422
rect 2741 418 2742 422
rect 2933 418 2934 422
rect 2994 418 2995 422
rect 3314 418 3315 422
rect 344 403 346 407
rect 350 403 353 407
rect 357 403 360 407
rect 1360 403 1362 407
rect 1366 403 1369 407
rect 1373 403 1376 407
rect 2384 403 2386 407
rect 2390 403 2393 407
rect 2397 403 2400 407
rect 3408 403 3410 407
rect 3414 403 3417 407
rect 3421 403 3424 407
rect 261 388 262 392
rect 3730 388 3732 392
rect 1022 371 1025 381
rect 1006 368 1025 371
rect 1146 368 1147 372
rect 1874 368 1875 372
rect 2090 368 2097 371
rect 2757 368 2758 372
rect 3349 368 3350 372
rect 1166 366 1170 368
rect 239 348 257 351
rect 830 348 846 351
rect 854 348 862 351
rect 874 348 894 351
rect 1046 351 1049 358
rect 1046 348 1057 351
rect 1126 348 1134 351
rect 1158 351 1161 361
rect 1578 358 1585 361
rect 1842 358 1849 361
rect 1886 358 1894 361
rect 2450 358 2454 362
rect 1158 348 1177 351
rect 1214 348 1222 351
rect 1282 348 1289 351
rect 1434 348 1446 351
rect 1890 348 1913 351
rect 2054 348 2062 351
rect 2158 348 2169 351
rect 2326 348 2334 351
rect 2358 348 2385 351
rect 2402 348 2425 351
rect 2454 348 2462 351
rect 2770 348 2785 351
rect 2846 351 2849 361
rect 2806 348 2833 351
rect 2846 348 2865 351
rect 2870 348 2878 351
rect 3246 351 3249 361
rect 3206 348 3233 351
rect 3246 348 3265 351
rect 3366 351 3369 358
rect 3358 348 3369 351
rect 3394 348 3401 351
rect 3450 348 3457 351
rect 3462 348 3470 351
rect 3614 348 3622 351
rect 882 338 889 341
rect 1182 338 1190 341
rect 1250 338 1265 341
rect 1342 338 1385 341
rect 1614 338 1633 341
rect 1954 338 1961 341
rect 2026 338 2033 341
rect 2150 338 2166 341
rect 2182 338 2201 341
rect 2222 338 2233 341
rect 2398 338 2414 341
rect 2462 338 2470 341
rect 2486 338 2502 341
rect 2914 338 2921 341
rect 3358 338 3361 348
rect 3414 338 3422 341
rect 3442 338 3449 341
rect 3662 338 3665 348
rect 270 328 286 331
rect 2118 328 2137 331
rect 1493 318 1494 322
rect 848 303 850 307
rect 854 303 857 307
rect 861 303 864 307
rect 1880 303 1882 307
rect 1886 303 1889 307
rect 1893 303 1896 307
rect 2904 303 2906 307
rect 2910 303 2913 307
rect 2917 303 2920 307
rect 1938 288 1939 292
rect 2021 288 2022 292
rect 3346 278 3369 281
rect 682 268 689 271
rect 1142 268 1153 271
rect 1606 268 1614 271
rect 2166 268 2185 271
rect 2799 268 2817 271
rect 2934 268 2942 271
rect 422 258 425 268
rect 3022 262 3025 271
rect 670 258 694 261
rect 702 258 721 261
rect 962 258 969 261
rect 1142 258 1150 261
rect 2046 258 2057 261
rect 2142 258 2153 261
rect 2174 258 2182 261
rect 2966 258 2985 261
rect 3046 261 3049 271
rect 3046 258 3065 261
rect 1182 248 1193 251
rect 1854 248 1865 251
rect 1918 248 1929 251
rect 2078 248 2089 251
rect 2098 248 2102 252
rect 2842 248 2846 252
rect 2898 248 2913 251
rect 1182 242 1185 248
rect 1862 242 1866 244
rect 1926 242 1929 248
rect 1026 238 1027 242
rect 1094 238 1113 241
rect 1890 238 1913 241
rect 1994 238 2001 241
rect 1110 228 1113 238
rect 562 218 563 222
rect 669 218 670 222
rect 1082 218 1083 222
rect 2258 218 2259 222
rect 2874 218 2875 222
rect 3005 218 3006 222
rect 3082 218 3083 222
rect 3290 218 3291 222
rect 344 203 346 207
rect 350 203 353 207
rect 357 203 360 207
rect 1360 203 1362 207
rect 1366 203 1369 207
rect 1373 203 1376 207
rect 2384 203 2386 207
rect 2390 203 2393 207
rect 2397 203 2400 207
rect 3408 203 3410 207
rect 3414 203 3417 207
rect 3421 203 3424 207
rect 1102 171 1105 181
rect 1102 168 1122 171
rect 1133 168 1134 172
rect 1658 168 1665 171
rect 618 158 622 162
rect 986 158 990 162
rect 1066 158 1070 162
rect 1214 152 1217 161
rect 602 148 617 151
rect 654 148 673 151
rect 730 148 737 151
rect 742 148 761 151
rect 1002 148 1009 151
rect 1134 148 1153 151
rect 1182 148 1190 151
rect 1250 148 1257 151
rect 1422 142 1425 151
rect 1814 148 1817 158
rect 2126 151 2129 161
rect 2210 158 2217 161
rect 2110 148 2129 151
rect 2694 148 2713 151
rect 2870 148 2878 151
rect 2962 148 2969 151
rect 3006 148 3014 151
rect 346 138 361 141
rect 1150 138 1169 141
rect 1226 138 1233 141
rect 2182 138 2185 148
rect 2846 141 2849 148
rect 2926 141 2929 148
rect 2846 138 2857 141
rect 2894 138 2929 141
rect 3314 138 3329 141
rect 3610 138 3617 141
rect 1014 128 1017 138
rect 2654 128 2673 131
rect 774 118 782 121
rect 848 103 850 107
rect 854 103 857 107
rect 861 103 864 107
rect 1880 103 1882 107
rect 1886 103 1889 107
rect 1893 103 1896 107
rect 2904 103 2906 107
rect 2910 103 2913 107
rect 2917 103 2920 107
rect 276 88 278 92
rect 2197 88 2198 92
rect 3326 88 3334 91
rect 3458 88 3460 92
rect 1998 78 2006 81
rect 2846 78 2854 81
rect 22 58 41 61
rect 246 61 249 71
rect 2878 71 2881 81
rect 2862 68 2881 71
rect 3566 68 3574 71
rect 246 58 258 61
rect 390 58 409 61
rect 999 58 1017 61
rect 1158 58 1161 68
rect 1199 58 1217 61
rect 1399 58 1433 61
rect 1711 58 1729 61
rect 2134 58 2137 68
rect 2630 58 2633 68
rect 3546 58 3553 61
rect 3730 58 3745 61
rect 254 56 258 58
rect 3354 48 3361 51
rect 344 3 346 7
rect 350 3 353 7
rect 357 3 360 7
rect 1360 3 1362 7
rect 1366 3 1369 7
rect 1373 3 1376 7
rect 2384 3 2386 7
rect 2390 3 2393 7
rect 2397 3 2400 7
rect 3408 3 3410 7
rect 3414 3 3417 7
rect 3421 3 3424 7
<< m2contact >>
rect 346 3603 350 3607
rect 353 3603 357 3607
rect 1362 3603 1366 3607
rect 1369 3603 1373 3607
rect 2386 3603 2390 3607
rect 2393 3603 2397 3607
rect 3410 3603 3414 3607
rect 3417 3603 3421 3607
rect 150 3588 154 3592
rect 262 3588 266 3592
rect 270 3588 274 3592
rect 294 3588 298 3592
rect 318 3588 322 3592
rect 534 3588 538 3592
rect 750 3588 754 3592
rect 758 3588 762 3592
rect 990 3588 994 3592
rect 1014 3588 1018 3592
rect 1190 3588 1194 3592
rect 1214 3588 1218 3592
rect 1238 3588 1242 3592
rect 1430 3588 1434 3592
rect 1454 3588 1458 3592
rect 1478 3588 1482 3592
rect 1502 3588 1506 3592
rect 1702 3588 1706 3592
rect 1726 3588 1730 3592
rect 1750 3588 1754 3592
rect 1942 3588 1946 3592
rect 1950 3588 1954 3592
rect 2702 3588 2706 3592
rect 3118 3588 3122 3592
rect 494 3579 498 3583
rect 694 3579 698 3583
rect 934 3579 938 3583
rect 1542 3579 1546 3583
rect 2230 3579 2234 3583
rect 2542 3579 2546 3583
rect 2990 3579 2994 3583
rect 3342 3578 3346 3582
rect 2446 3568 2450 3572
rect 3198 3568 3202 3572
rect 3230 3568 3234 3572
rect 3486 3568 3490 3572
rect 3670 3568 3674 3572
rect 494 3556 498 3560
rect 694 3556 698 3560
rect 934 3556 938 3560
rect 1014 3558 1018 3562
rect 1238 3558 1242 3562
rect 1542 3556 1546 3560
rect 1750 3558 1754 3562
rect 2230 3556 2234 3560
rect 2374 3558 2378 3562
rect 2398 3558 2402 3562
rect 2462 3558 2466 3562
rect 2478 3558 2482 3562
rect 2542 3556 2546 3560
rect 2702 3558 2706 3562
rect 2902 3558 2906 3562
rect 166 3548 170 3552
rect 174 3548 178 3552
rect 246 3548 250 3552
rect 286 3548 290 3552
rect 310 3548 314 3552
rect 510 3548 514 3552
rect 606 3548 610 3552
rect 734 3548 738 3552
rect 942 3548 946 3552
rect 974 3548 978 3552
rect 1014 3548 1018 3552
rect 1118 3548 1122 3552
rect 1159 3548 1163 3552
rect 1166 3548 1170 3552
rect 1198 3548 1202 3552
rect 1238 3548 1242 3552
rect 1342 3548 1346 3552
rect 1383 3548 1387 3552
rect 1398 3548 1402 3552
rect 1438 3548 1442 3552
rect 1462 3548 1466 3552
rect 1486 3548 1490 3552
rect 1526 3548 1530 3552
rect 1630 3548 1634 3552
rect 1710 3548 1714 3552
rect 1750 3548 1754 3552
rect 1966 3548 1970 3552
rect 1998 3548 2002 3552
rect 2190 3548 2194 3552
rect 2222 3548 2226 3552
rect 2430 3548 2434 3552
rect 2446 3548 2450 3552
rect 2462 3548 2466 3552
rect 2502 3548 2506 3552
rect 2630 3548 2634 3552
rect 2702 3548 2706 3552
rect 2806 3548 2810 3552
rect 2862 3548 2866 3552
rect 2886 3548 2890 3552
rect 2990 3556 2994 3560
rect 3158 3558 3162 3562
rect 3182 3558 3186 3562
rect 2942 3548 2946 3552
rect 2974 3548 2978 3552
rect 3150 3548 3154 3552
rect 3198 3548 3202 3552
rect 3278 3558 3282 3562
rect 3318 3558 3322 3562
rect 3334 3558 3338 3562
rect 3390 3558 3394 3562
rect 3470 3558 3474 3562
rect 3654 3558 3658 3562
rect 3230 3548 3234 3552
rect 3262 3548 3266 3552
rect 3358 3548 3362 3552
rect 3422 3548 3426 3552
rect 3462 3548 3466 3552
rect 3478 3548 3482 3552
rect 3502 3548 3506 3552
rect 3526 3548 3530 3552
rect 3550 3548 3554 3552
rect 3574 3548 3578 3552
rect 3614 3548 3618 3552
rect 3646 3548 3650 3552
rect 3662 3548 3666 3552
rect 3710 3548 3714 3552
rect 6 3538 10 3542
rect 70 3538 74 3542
rect 78 3538 82 3542
rect 238 3538 242 3542
rect 462 3538 466 3542
rect 662 3538 666 3542
rect 902 3538 906 3542
rect 1062 3538 1066 3542
rect 1286 3538 1290 3542
rect 1574 3538 1578 3542
rect 1798 3538 1802 3542
rect 1990 3538 1994 3542
rect 2022 3538 2026 3542
rect 2094 3538 2098 3542
rect 2166 3538 2170 3542
rect 2262 3538 2266 3542
rect 2390 3538 2394 3542
rect 2422 3538 2426 3542
rect 2438 3538 2442 3542
rect 2478 3538 2482 3542
rect 2494 3538 2498 3542
rect 2574 3538 2578 3542
rect 2750 3538 2754 3542
rect 2886 3538 2890 3542
rect 2910 3538 2914 3542
rect 2950 3538 2954 3542
rect 3022 3538 3026 3542
rect 3158 3538 3162 3542
rect 3174 3538 3178 3542
rect 3206 3538 3210 3542
rect 3246 3538 3250 3542
rect 3254 3538 3258 3542
rect 3286 3538 3290 3542
rect 3294 3538 3298 3542
rect 3318 3538 3322 3542
rect 3326 3538 3330 3542
rect 3366 3538 3370 3542
rect 3454 3538 3458 3542
rect 3542 3538 3546 3542
rect 3734 3540 3738 3544
rect 3742 3538 3746 3542
rect 446 3528 450 3532
rect 646 3528 650 3532
rect 886 3528 890 3532
rect 1078 3528 1082 3532
rect 1302 3528 1306 3532
rect 1590 3528 1594 3532
rect 1814 3528 1818 3532
rect 1974 3528 1978 3532
rect 2014 3528 2018 3532
rect 2174 3528 2178 3532
rect 2278 3528 2282 3532
rect 2590 3528 2594 3532
rect 2766 3528 2770 3532
rect 2862 3528 2866 3532
rect 3038 3528 3042 3532
rect 3150 3528 3154 3532
rect 3310 3528 3314 3532
rect 3414 3528 3418 3532
rect 3438 3528 3442 3532
rect 3446 3528 3450 3532
rect 3478 3528 3482 3532
rect 3518 3528 3522 3532
rect 3590 3528 3594 3532
rect 3598 3528 3602 3532
rect 134 3518 138 3522
rect 1982 3518 1986 3522
rect 2038 3518 2042 3522
rect 2182 3518 2186 3522
rect 2358 3518 2362 3522
rect 2670 3518 2674 3522
rect 2846 3518 2850 3522
rect 3118 3518 3122 3522
rect 3510 3518 3514 3522
rect 3566 3518 3570 3522
rect 3582 3518 3586 3522
rect 3606 3518 3610 3522
rect 3630 3518 3634 3522
rect 3670 3518 3674 3522
rect 3694 3518 3698 3522
rect 3718 3518 3722 3522
rect 850 3503 854 3507
rect 857 3503 861 3507
rect 1882 3503 1886 3507
rect 1889 3503 1893 3507
rect 2906 3503 2910 3507
rect 2913 3503 2917 3507
rect 206 3488 210 3492
rect 422 3488 426 3492
rect 1166 3488 1170 3492
rect 1230 3488 1234 3492
rect 1270 3488 1274 3492
rect 1302 3488 1306 3492
rect 1350 3488 1354 3492
rect 2230 3488 2234 3492
rect 2246 3488 2250 3492
rect 2278 3488 2282 3492
rect 2830 3488 2834 3492
rect 2862 3488 2866 3492
rect 2926 3488 2930 3492
rect 3646 3488 3650 3492
rect 3686 3488 3690 3492
rect 318 3478 322 3482
rect 534 3478 538 3482
rect 702 3478 706 3482
rect 894 3478 898 3482
rect 1070 3478 1074 3482
rect 1238 3478 1242 3482
rect 1438 3478 1442 3482
rect 1614 3478 1618 3482
rect 1710 3478 1714 3482
rect 1798 3478 1802 3482
rect 1990 3478 1994 3482
rect 2182 3478 2186 3482
rect 2238 3478 2242 3482
rect 2270 3478 2274 3482
rect 2302 3478 2306 3482
rect 2350 3478 2354 3482
rect 2438 3478 2442 3482
rect 2526 3478 2530 3482
rect 2662 3478 2666 3482
rect 2902 3478 2906 3482
rect 3078 3478 3082 3482
rect 3150 3478 3154 3482
rect 3158 3478 3162 3482
rect 30 3468 34 3472
rect 102 3468 106 3472
rect 166 3468 170 3472
rect 334 3468 338 3472
rect 550 3468 554 3472
rect 686 3468 690 3472
rect 878 3468 882 3472
rect 1054 3468 1058 3472
rect 1214 3468 1218 3472
rect 1246 3468 1250 3472
rect 1278 3468 1282 3472
rect 1310 3468 1314 3472
rect 1422 3468 1426 3472
rect 1478 3468 1482 3472
rect 1598 3468 1602 3472
rect 1814 3468 1818 3472
rect 2006 3468 2010 3472
rect 2142 3468 2146 3472
rect 2206 3468 2210 3472
rect 2254 3468 2258 3472
rect 2262 3468 2266 3472
rect 2454 3468 2458 3472
rect 2534 3468 2538 3472
rect 2574 3468 2578 3472
rect 2646 3468 2650 3472
rect 2790 3468 2794 3472
rect 2854 3468 2858 3472
rect 2878 3468 2882 3472
rect 2950 3468 2954 3472
rect 3014 3468 3018 3472
rect 3062 3468 3066 3472
rect 3118 3468 3122 3472
rect 3142 3468 3146 3472
rect 22 3458 26 3462
rect 198 3458 202 3462
rect 382 3458 386 3462
rect 438 3458 442 3462
rect 582 3458 586 3462
rect 598 3458 602 3462
rect 366 3450 370 3454
rect 742 3458 746 3462
rect 846 3458 850 3462
rect 934 3458 938 3462
rect 1014 3458 1018 3462
rect 1110 3458 1114 3462
rect 1206 3458 1210 3462
rect 1222 3458 1226 3462
rect 1238 3458 1242 3462
rect 1254 3458 1258 3462
rect 1286 3458 1290 3462
rect 1318 3458 1322 3462
rect 1374 3458 1378 3462
rect 1550 3458 1554 3462
rect 1862 3458 1866 3462
rect 2046 3458 2050 3462
rect 2150 3458 2154 3462
rect 2198 3458 2202 3462
rect 2214 3458 2218 3462
rect 2262 3458 2266 3462
rect 2486 3458 2490 3462
rect 2542 3458 2546 3462
rect 2550 3458 2554 3462
rect 2566 3458 2570 3462
rect 2606 3458 2610 3462
rect 2702 3458 2706 3462
rect 2758 3458 2762 3462
rect 2798 3458 2802 3462
rect 2830 3458 2834 3462
rect 2846 3458 2850 3462
rect 2886 3458 2890 3462
rect 2998 3458 3002 3462
rect 3006 3458 3010 3462
rect 3062 3458 3066 3462
rect 3078 3458 3082 3462
rect 3118 3458 3122 3462
rect 3174 3458 3178 3462
rect 3190 3458 3194 3462
rect 3230 3458 3234 3462
rect 3254 3458 3258 3462
rect 3294 3458 3298 3462
rect 3310 3468 3314 3472
rect 3382 3468 3386 3472
rect 3390 3468 3394 3472
rect 3430 3478 3434 3482
rect 3510 3478 3514 3482
rect 3726 3478 3730 3482
rect 3438 3468 3442 3472
rect 3462 3468 3466 3472
rect 3518 3468 3522 3472
rect 3622 3468 3626 3472
rect 3662 3468 3666 3472
rect 3742 3468 3746 3472
rect 3758 3468 3762 3472
rect 3310 3458 3314 3462
rect 3326 3458 3330 3462
rect 3350 3458 3354 3462
rect 3478 3458 3482 3462
rect 3542 3458 3546 3462
rect 3566 3458 3570 3462
rect 3606 3458 3610 3462
rect 3670 3458 3674 3462
rect 3702 3458 3706 3462
rect 3750 3458 3754 3462
rect 598 3448 602 3452
rect 630 3448 634 3452
rect 638 3448 642 3452
rect 830 3448 834 3452
rect 1022 3450 1026 3454
rect 1190 3448 1194 3452
rect 1270 3448 1274 3452
rect 1302 3448 1306 3452
rect 1334 3448 1338 3452
rect 1390 3450 1394 3454
rect 1566 3450 1570 3454
rect 1846 3450 1850 3454
rect 2054 3448 2058 3452
rect 2502 3448 2506 3452
rect 2550 3448 2554 3452
rect 2598 3448 2602 3452
rect 2814 3448 2818 3452
rect 2862 3448 2866 3452
rect 2934 3448 2938 3452
rect 2958 3448 2962 3452
rect 2982 3448 2986 3452
rect 3014 3448 3018 3452
rect 3038 3448 3042 3452
rect 3126 3448 3130 3452
rect 3206 3448 3210 3452
rect 3222 3448 3226 3452
rect 3270 3448 3274 3452
rect 3278 3448 3282 3452
rect 3326 3448 3330 3452
rect 3358 3448 3362 3452
rect 3494 3448 3498 3452
rect 3542 3448 3546 3452
rect 3582 3448 3586 3452
rect 3614 3448 3618 3452
rect 3686 3448 3690 3452
rect 3694 3448 3698 3452
rect 3774 3448 3778 3452
rect 6 3438 10 3442
rect 982 3438 986 3442
rect 2166 3438 2170 3442
rect 3230 3438 3234 3442
rect 3262 3438 3266 3442
rect 3342 3438 3346 3442
rect 3534 3438 3538 3442
rect 3566 3438 3570 3442
rect 3590 3438 3594 3442
rect 3598 3438 3602 3442
rect 3710 3438 3714 3442
rect 366 3427 370 3431
rect 1022 3427 1026 3431
rect 1150 3428 1154 3432
rect 1390 3427 1394 3431
rect 1518 3428 1522 3432
rect 2742 3428 2746 3432
rect 86 3418 90 3422
rect 182 3418 186 3422
rect 454 3418 458 3422
rect 598 3418 602 3422
rect 638 3418 642 3422
rect 782 3418 786 3422
rect 830 3418 834 3422
rect 1566 3418 1570 3422
rect 1718 3418 1722 3422
rect 1846 3418 1850 3422
rect 1910 3418 1914 3422
rect 2054 3418 2058 3422
rect 2086 3418 2090 3422
rect 2310 3418 2314 3422
rect 2358 3418 2362 3422
rect 2502 3418 2506 3422
rect 2598 3418 2602 3422
rect 2774 3418 2778 3422
rect 2966 3418 2970 3422
rect 3022 3418 3026 3422
rect 3190 3418 3194 3422
rect 3238 3418 3242 3422
rect 3262 3418 3266 3422
rect 3294 3418 3298 3422
rect 3350 3418 3354 3422
rect 3398 3418 3402 3422
rect 3454 3418 3458 3422
rect 3486 3418 3490 3422
rect 3542 3418 3546 3422
rect 3574 3418 3578 3422
rect 3630 3418 3634 3422
rect 3702 3418 3706 3422
rect 3726 3418 3730 3422
rect 3766 3418 3770 3422
rect 346 3403 350 3407
rect 353 3403 357 3407
rect 1362 3403 1366 3407
rect 1369 3403 1373 3407
rect 2386 3403 2390 3407
rect 2393 3403 2397 3407
rect 3410 3403 3414 3407
rect 3417 3403 3421 3407
rect 222 3388 226 3392
rect 294 3388 298 3392
rect 326 3388 330 3392
rect 374 3388 378 3392
rect 406 3388 410 3392
rect 646 3388 650 3392
rect 670 3388 674 3392
rect 1014 3388 1018 3392
rect 1062 3388 1066 3392
rect 1094 3388 1098 3392
rect 1238 3388 1242 3392
rect 1270 3388 1274 3392
rect 1398 3388 1402 3392
rect 1542 3388 1546 3392
rect 1582 3388 1586 3392
rect 1742 3388 1746 3392
rect 1950 3388 1954 3392
rect 2190 3388 2194 3392
rect 2590 3388 2594 3392
rect 2950 3388 2954 3392
rect 566 3379 570 3383
rect 830 3379 834 3383
rect 6 3368 10 3372
rect 30 3368 34 3372
rect 926 3368 930 3372
rect 1622 3378 1626 3382
rect 1822 3379 1826 3383
rect 2142 3379 2146 3383
rect 2342 3379 2346 3383
rect 2646 3379 2650 3383
rect 3318 3378 3322 3382
rect 1310 3368 1314 3372
rect 1606 3368 1610 3372
rect 2782 3368 2786 3372
rect 3102 3368 3106 3372
rect 3206 3368 3210 3372
rect 3214 3368 3218 3372
rect 3262 3368 3266 3372
rect 3310 3368 3314 3372
rect 3430 3368 3434 3372
rect 3742 3368 3746 3372
rect 222 3358 226 3362
rect 310 3358 314 3362
rect 342 3358 346 3362
rect 390 3358 394 3362
rect 566 3356 570 3360
rect 606 3358 610 3362
rect 630 3358 634 3362
rect 830 3356 834 3360
rect 942 3358 946 3362
rect 1054 3358 1058 3362
rect 1238 3358 1242 3362
rect 1294 3358 1298 3362
rect 1366 3358 1370 3362
rect 1542 3358 1546 3362
rect 1590 3358 1594 3362
rect 1822 3356 1826 3360
rect 1974 3358 1978 3362
rect 1990 3358 1994 3362
rect 2142 3356 2146 3360
rect 2342 3356 2346 3360
rect 2398 3358 2402 3362
rect 2590 3358 2594 3362
rect 2646 3356 2650 3360
rect 3006 3358 3010 3362
rect 3118 3358 3122 3362
rect 3126 3358 3130 3362
rect 3222 3358 3226 3362
rect 3246 3358 3250 3362
rect 3278 3358 3282 3362
rect 3294 3358 3298 3362
rect 3374 3358 3378 3362
rect 3406 3358 3410 3362
rect 3430 3358 3434 3362
rect 3478 3358 3482 3362
rect 3526 3358 3530 3362
rect 3566 3358 3570 3362
rect 3726 3358 3730 3362
rect 3750 3358 3754 3362
rect 22 3348 26 3352
rect 54 3348 58 3352
rect 206 3348 210 3352
rect 254 3348 258 3352
rect 270 3348 274 3352
rect 286 3348 290 3352
rect 318 3348 322 3352
rect 374 3348 378 3352
rect 422 3348 426 3352
rect 582 3348 586 3352
rect 646 3348 650 3352
rect 742 3348 746 3352
rect 846 3348 850 3352
rect 886 3348 890 3352
rect 934 3348 938 3352
rect 998 3348 1002 3352
rect 1038 3348 1042 3352
rect 1054 3348 1058 3352
rect 1086 3348 1090 3352
rect 1134 3348 1138 3352
rect 1270 3348 1274 3352
rect 1302 3348 1306 3352
rect 1326 3348 1330 3352
rect 1350 3348 1354 3352
rect 1366 3348 1370 3352
rect 1526 3348 1530 3352
rect 1566 3348 1570 3352
rect 1758 3348 1762 3352
rect 1806 3348 1810 3352
rect 2054 3348 2058 3352
rect 2150 3348 2154 3352
rect 2182 3348 2186 3352
rect 2254 3348 2258 3352
rect 2358 3348 2362 3352
rect 2486 3348 2490 3352
rect 2590 3348 2594 3352
rect 2638 3348 2642 3352
rect 2734 3348 2738 3352
rect 2870 3348 2874 3352
rect 2878 3348 2882 3352
rect 2886 3348 2890 3352
rect 2918 3348 2922 3352
rect 2950 3348 2954 3352
rect 2966 3348 2970 3352
rect 2998 3348 3002 3352
rect 3022 3348 3026 3352
rect 3110 3348 3114 3352
rect 3174 3348 3178 3352
rect 3214 3348 3218 3352
rect 3270 3348 3274 3352
rect 3318 3348 3322 3352
rect 3358 3348 3362 3352
rect 3382 3348 3386 3352
rect 3438 3348 3442 3352
rect 3558 3348 3562 3352
rect 3598 3348 3602 3352
rect 3622 3348 3626 3352
rect 3670 3348 3674 3352
rect 3678 3348 3682 3352
rect 3758 3348 3762 3352
rect 77 3338 81 3342
rect 174 3338 178 3342
rect 246 3338 250 3342
rect 278 3338 282 3342
rect 286 3338 290 3342
rect 318 3338 322 3342
rect 366 3338 370 3342
rect 534 3338 538 3342
rect 622 3338 626 3342
rect 654 3338 658 3342
rect 798 3338 802 3342
rect 958 3338 962 3342
rect 974 3338 978 3342
rect 982 3338 986 3342
rect 1030 3338 1034 3342
rect 1190 3338 1194 3342
rect 1262 3338 1266 3342
rect 1494 3338 1498 3342
rect 1590 3338 1594 3342
rect 1678 3338 1682 3342
rect 1782 3338 1786 3342
rect 1854 3338 1858 3342
rect 1998 3338 2002 3342
rect 2110 3338 2114 3342
rect 2310 3338 2314 3342
rect 2382 3338 2386 3342
rect 2542 3338 2546 3342
rect 2678 3338 2682 3342
rect 2790 3338 2794 3342
rect 2854 3338 2858 3342
rect 2862 3338 2866 3342
rect 2894 3338 2898 3342
rect 2910 3338 2914 3342
rect 2942 3338 2946 3342
rect 3030 3338 3034 3342
rect 3086 3338 3090 3342
rect 3142 3338 3146 3342
rect 3166 3338 3170 3342
rect 3190 3338 3194 3342
rect 3230 3338 3234 3342
rect 3270 3338 3274 3342
rect 3334 3338 3338 3342
rect 3342 3338 3346 3342
rect 3350 3338 3354 3342
rect 3382 3338 3386 3342
rect 3462 3338 3466 3342
rect 3486 3338 3490 3342
rect 3510 3338 3514 3342
rect 3526 3338 3530 3342
rect 3550 3338 3554 3342
rect 3582 3338 3586 3342
rect 3590 3338 3594 3342
rect 3630 3338 3634 3342
rect 3686 3338 3690 3342
rect 3718 3338 3722 3342
rect 3742 3338 3746 3342
rect 3758 3338 3762 3342
rect 54 3328 58 3332
rect 70 3328 74 3332
rect 158 3328 162 3332
rect 438 3328 442 3332
rect 518 3328 522 3332
rect 782 3328 786 3332
rect 982 3328 986 3332
rect 1174 3328 1178 3332
rect 1326 3328 1330 3332
rect 1478 3328 1482 3332
rect 1870 3328 1874 3332
rect 2094 3328 2098 3332
rect 2198 3328 2202 3332
rect 2294 3328 2298 3332
rect 2438 3328 2442 3332
rect 2526 3328 2530 3332
rect 2694 3328 2698 3332
rect 2934 3328 2938 3332
rect 2982 3328 2986 3332
rect 2998 3328 3002 3332
rect 3150 3328 3154 3332
rect 3294 3328 3298 3332
rect 3486 3328 3490 3332
rect 3534 3328 3538 3332
rect 3646 3328 3650 3332
rect 3654 3328 3658 3332
rect 3710 3328 3714 3332
rect 270 3318 274 3322
rect 606 3318 610 3322
rect 702 3318 706 3322
rect 902 3318 906 3322
rect 1398 3318 1402 3322
rect 2014 3318 2018 3322
rect 2214 3318 2218 3322
rect 2390 3318 2394 3322
rect 2414 3318 2418 3322
rect 2446 3318 2450 3322
rect 3054 3318 3058 3322
rect 3094 3318 3098 3322
rect 3182 3318 3186 3322
rect 3206 3318 3210 3322
rect 3374 3318 3378 3322
rect 3406 3318 3410 3322
rect 3446 3318 3450 3322
rect 3542 3318 3546 3322
rect 3566 3318 3570 3322
rect 3614 3318 3618 3322
rect 3638 3318 3642 3322
rect 3662 3318 3666 3322
rect 3694 3318 3698 3322
rect 3726 3318 3730 3322
rect 850 3303 854 3307
rect 857 3303 861 3307
rect 1882 3303 1886 3307
rect 1889 3303 1893 3307
rect 2906 3303 2910 3307
rect 2913 3303 2917 3307
rect 222 3288 226 3292
rect 398 3288 402 3292
rect 414 3288 418 3292
rect 454 3288 458 3292
rect 662 3288 666 3292
rect 862 3288 866 3292
rect 1190 3288 1194 3292
rect 1230 3288 1234 3292
rect 1374 3288 1378 3292
rect 1422 3288 1426 3292
rect 1510 3288 1514 3292
rect 2494 3288 2498 3292
rect 2622 3288 2626 3292
rect 2638 3288 2642 3292
rect 2678 3288 2682 3292
rect 2902 3288 2906 3292
rect 2950 3288 2954 3292
rect 2974 3288 2978 3292
rect 3014 3288 3018 3292
rect 3318 3288 3322 3292
rect 3742 3288 3746 3292
rect 118 3278 122 3282
rect 318 3278 322 3282
rect 534 3278 538 3282
rect 942 3278 946 3282
rect 1110 3278 1114 3282
rect 1238 3278 1242 3282
rect 1462 3278 1466 3282
rect 1790 3278 1794 3282
rect 2006 3278 2010 3282
rect 2182 3278 2186 3282
rect 2334 3278 2338 3282
rect 2350 3278 2354 3282
rect 2398 3278 2402 3282
rect 2446 3278 2450 3282
rect 2510 3278 2514 3282
rect 2526 3278 2530 3282
rect 2574 3278 2578 3282
rect 2782 3278 2786 3282
rect 2990 3278 2994 3282
rect 3006 3278 3010 3282
rect 3310 3278 3314 3282
rect 3350 3278 3354 3282
rect 3470 3278 3474 3282
rect 3478 3278 3482 3282
rect 3502 3278 3506 3282
rect 3630 3278 3634 3282
rect 3638 3278 3642 3282
rect 3750 3278 3754 3282
rect 134 3268 138 3272
rect 302 3268 306 3272
rect 446 3268 450 3272
rect 478 3268 482 3272
rect 502 3268 506 3272
rect 518 3268 522 3272
rect 550 3268 554 3272
rect 582 3268 586 3272
rect 598 3268 602 3272
rect 614 3268 618 3272
rect 654 3268 658 3272
rect 686 3268 690 3272
rect 694 3268 698 3272
rect 710 3268 714 3272
rect 774 3268 778 3272
rect 782 3268 786 3272
rect 798 3268 802 3272
rect 814 3268 818 3272
rect 830 3268 834 3272
rect 958 3268 962 3272
rect 1094 3268 1098 3272
rect 1206 3268 1210 3272
rect 1286 3268 1290 3272
rect 1302 3268 1306 3272
rect 1318 3268 1322 3272
rect 1342 3268 1346 3272
rect 1446 3268 1450 3272
rect 1486 3268 1490 3272
rect 1606 3268 1610 3272
rect 1670 3268 1674 3272
rect 1806 3268 1810 3272
rect 1910 3268 1914 3272
rect 2022 3268 2026 3272
rect 2198 3268 2202 3272
rect 2294 3268 2298 3272
rect 2302 3268 2306 3272
rect 2318 3268 2322 3272
rect 2374 3268 2378 3272
rect 2414 3268 2418 3272
rect 2446 3268 2450 3272
rect 2518 3268 2522 3272
rect 2798 3268 2802 3272
rect 2870 3268 2874 3272
rect 2918 3268 2922 3272
rect 2958 3268 2962 3272
rect 2966 3268 2970 3272
rect 3038 3268 3042 3272
rect 3046 3268 3050 3272
rect 3086 3268 3090 3272
rect 3118 3268 3122 3272
rect 3126 3268 3130 3272
rect 3182 3268 3186 3272
rect 3206 3268 3210 3272
rect 3222 3268 3226 3272
rect 3286 3268 3290 3272
rect 3294 3268 3298 3272
rect 3334 3266 3338 3270
rect 3342 3268 3346 3272
rect 3406 3268 3410 3272
rect 3518 3268 3522 3272
rect 3646 3268 3650 3272
rect 3686 3268 3690 3272
rect 3734 3268 3738 3272
rect 174 3258 178 3262
rect 206 3258 210 3262
rect 358 3258 362 3262
rect 470 3258 474 3262
rect 614 3258 618 3262
rect 630 3258 634 3262
rect 678 3258 682 3262
rect 718 3258 722 3262
rect 758 3258 762 3262
rect 806 3258 810 3262
rect 830 3258 834 3262
rect 902 3258 906 3262
rect 1046 3258 1050 3262
rect 1214 3258 1218 3262
rect 1238 3258 1242 3262
rect 1262 3258 1266 3262
rect 1294 3258 1298 3262
rect 1350 3258 1354 3262
rect 1406 3258 1410 3262
rect 1478 3258 1482 3262
rect 1526 3258 1530 3262
rect 1630 3258 1634 3262
rect 1638 3258 1642 3262
rect 1662 3258 1666 3262
rect 1694 3258 1698 3262
rect 1846 3258 1850 3262
rect 2054 3258 2058 3262
rect 2142 3258 2146 3262
rect 2254 3258 2258 3262
rect 2294 3258 2298 3262
rect 2310 3258 2314 3262
rect 2350 3258 2354 3262
rect 2366 3258 2370 3262
rect 2422 3258 2426 3262
rect 2470 3258 2474 3262
rect 2478 3258 2482 3262
rect 2550 3258 2554 3262
rect 2566 3258 2570 3262
rect 2590 3258 2594 3262
rect 2598 3258 2602 3262
rect 2654 3258 2658 3262
rect 2742 3258 2746 3262
rect 2990 3258 2994 3262
rect 3030 3258 3034 3262
rect 3062 3258 3066 3262
rect 3102 3258 3106 3262
rect 3110 3258 3114 3262
rect 3158 3258 3162 3262
rect 3182 3258 3186 3262
rect 3238 3258 3242 3262
rect 3278 3258 3282 3262
rect 3294 3258 3298 3262
rect 3374 3258 3378 3262
rect 3430 3258 3434 3262
rect 3454 3258 3458 3262
rect 3470 3258 3474 3262
rect 3494 3258 3498 3262
rect 3526 3258 3530 3262
rect 3542 3258 3546 3262
rect 3582 3258 3586 3262
rect 3614 3258 3618 3262
rect 3654 3258 3658 3262
rect 3678 3258 3682 3262
rect 3710 3258 3714 3262
rect 3726 3258 3730 3262
rect 3774 3258 3778 3262
rect 182 3248 186 3252
rect 270 3250 274 3254
rect 430 3248 434 3252
rect 454 3248 458 3252
rect 510 3248 514 3252
rect 574 3248 578 3252
rect 606 3248 610 3252
rect 662 3248 666 3252
rect 766 3248 770 3252
rect 790 3248 794 3252
rect 990 3250 994 3254
rect 1014 3248 1018 3252
rect 1062 3250 1066 3254
rect 1230 3248 1234 3252
rect 1254 3248 1258 3252
rect 1334 3248 1338 3252
rect 1366 3248 1370 3252
rect 1414 3248 1418 3252
rect 1494 3248 1498 3252
rect 1542 3248 1546 3252
rect 1838 3250 1842 3254
rect 1894 3248 1898 3252
rect 2070 3248 2074 3252
rect 2230 3250 2234 3254
rect 2270 3248 2274 3252
rect 2286 3248 2290 3252
rect 2326 3248 2330 3252
rect 2390 3248 2394 3252
rect 2438 3248 2442 3252
rect 2494 3248 2498 3252
rect 2502 3248 2506 3252
rect 2566 3248 2570 3252
rect 2622 3248 2626 3252
rect 2830 3250 2834 3254
rect 3014 3248 3018 3252
rect 3094 3248 3098 3252
rect 3126 3248 3130 3252
rect 3142 3248 3146 3252
rect 3174 3248 3178 3252
rect 3198 3248 3202 3252
rect 3222 3248 3226 3252
rect 3238 3248 3242 3252
rect 3262 3248 3266 3252
rect 3382 3248 3386 3252
rect 3398 3248 3402 3252
rect 3534 3248 3538 3252
rect 3590 3248 3594 3252
rect 3606 3248 3610 3252
rect 3622 3248 3626 3252
rect 3662 3248 3666 3252
rect 3718 3248 3722 3252
rect 3766 3248 3770 3252
rect 6 3238 10 3242
rect 534 3238 538 3242
rect 750 3238 754 3242
rect 1262 3238 1266 3242
rect 1270 3238 1274 3242
rect 1398 3238 1402 3242
rect 3438 3238 3442 3242
rect 3550 3238 3554 3242
rect 3574 3238 3578 3242
rect 3614 3238 3618 3242
rect 270 3227 274 3231
rect 718 3228 722 3232
rect 990 3227 994 3231
rect 1062 3227 1066 3231
rect 2230 3227 2234 3231
rect 3542 3228 3546 3232
rect 182 3218 186 3222
rect 702 3218 706 3222
rect 1190 3218 1194 3222
rect 1614 3218 1618 3222
rect 1646 3218 1650 3222
rect 1710 3218 1714 3222
rect 1838 3218 1842 3222
rect 1902 3218 1906 3222
rect 1926 3218 1930 3222
rect 2070 3218 2074 3222
rect 2102 3218 2106 3222
rect 2702 3218 2706 3222
rect 2830 3218 2834 3222
rect 3054 3218 3058 3222
rect 3158 3218 3162 3222
rect 3214 3218 3218 3222
rect 3318 3218 3322 3222
rect 3350 3218 3354 3222
rect 3430 3218 3434 3222
rect 3486 3218 3490 3222
rect 3502 3218 3506 3222
rect 3582 3218 3586 3222
rect 3598 3218 3602 3222
rect 3678 3218 3682 3222
rect 3750 3218 3754 3222
rect 346 3203 350 3207
rect 353 3203 357 3207
rect 1362 3203 1366 3207
rect 1369 3203 1373 3207
rect 2386 3203 2390 3207
rect 2393 3203 2397 3207
rect 3410 3203 3414 3207
rect 3417 3203 3421 3207
rect 134 3188 138 3192
rect 358 3188 362 3192
rect 534 3188 538 3192
rect 678 3188 682 3192
rect 774 3188 778 3192
rect 798 3188 802 3192
rect 1166 3188 1170 3192
rect 1214 3188 1218 3192
rect 1510 3188 1514 3192
rect 1606 3188 1610 3192
rect 1718 3188 1722 3192
rect 2038 3188 2042 3192
rect 2174 3188 2178 3192
rect 2294 3188 2298 3192
rect 2646 3188 2650 3192
rect 3230 3188 3234 3192
rect 3558 3188 3562 3192
rect 3718 3188 3722 3192
rect 182 3179 186 3183
rect 734 3168 738 3172
rect 750 3168 754 3172
rect 806 3168 810 3172
rect 1038 3179 1042 3183
rect 886 3168 890 3172
rect 918 3168 922 3172
rect 1382 3168 1386 3172
rect 2726 3179 2730 3183
rect 1454 3168 1458 3172
rect 1518 3168 1522 3172
rect 1542 3168 1546 3172
rect 1726 3168 1730 3172
rect 1814 3168 1818 3172
rect 2214 3168 2218 3172
rect 2326 3168 2330 3172
rect 2398 3168 2402 3172
rect 3262 3168 3266 3172
rect 3550 3168 3554 3172
rect 3718 3168 3722 3172
rect 3726 3168 3730 3172
rect 182 3156 186 3160
rect 358 3158 362 3162
rect 534 3158 538 3162
rect 750 3158 754 3162
rect 758 3158 762 3162
rect 790 3158 794 3162
rect 870 3158 874 3162
rect 982 3158 986 3162
rect 998 3158 1002 3162
rect 1038 3156 1042 3160
rect 1214 3158 1218 3162
rect 1438 3158 1442 3162
rect 1494 3158 1498 3162
rect 1502 3158 1506 3162
rect 1750 3158 1754 3162
rect 1790 3158 1794 3162
rect 1798 3158 1802 3162
rect 1862 3158 1866 3162
rect 174 3148 178 3152
rect 270 3148 274 3152
rect 366 3148 370 3152
rect 534 3148 538 3152
rect 702 3148 706 3152
rect 742 3148 746 3152
rect 774 3148 778 3152
rect 798 3148 802 3152
rect 830 3148 834 3152
rect 878 3148 882 3152
rect 966 3148 970 3152
rect 982 3148 986 3152
rect 1022 3148 1026 3152
rect 1214 3148 1218 3152
rect 1414 3148 1418 3152
rect 1430 3148 1434 3152
rect 1446 3148 1450 3152
rect 1478 3148 1482 3152
rect 1494 3148 1498 3152
rect 1646 3148 1650 3152
rect 1686 3148 1690 3152
rect 1710 3148 1714 3152
rect 1734 3148 1738 3152
rect 1846 3148 1850 3152
rect 1958 3158 1962 3162
rect 1886 3148 1890 3152
rect 1926 3148 1930 3152
rect 1998 3158 2002 3162
rect 2022 3158 2026 3162
rect 2070 3158 2074 3162
rect 2078 3158 2082 3162
rect 2110 3158 2114 3162
rect 2158 3158 2162 3162
rect 2190 3158 2194 3162
rect 2198 3158 2202 3162
rect 2230 3158 2234 3162
rect 2270 3158 2274 3162
rect 1982 3148 1986 3152
rect 2038 3148 2042 3152
rect 2078 3148 2082 3152
rect 2102 3148 2106 3152
rect 2142 3148 2146 3152
rect 2214 3148 2218 3152
rect 2342 3158 2346 3162
rect 2382 3158 2386 3162
rect 2414 3158 2418 3162
rect 2510 3158 2514 3162
rect 2566 3158 2570 3162
rect 2574 3158 2578 3162
rect 2606 3158 2610 3162
rect 2294 3148 2298 3152
rect 2374 3148 2378 3152
rect 2398 3148 2402 3152
rect 2438 3148 2442 3152
rect 2486 3148 2490 3152
rect 2510 3148 2514 3152
rect 2534 3148 2538 3152
rect 2550 3148 2554 3152
rect 2574 3148 2578 3152
rect 2622 3148 2626 3152
rect 2646 3148 2650 3152
rect 2670 3158 2674 3162
rect 2726 3156 2730 3160
rect 2926 3158 2930 3162
rect 3014 3158 3018 3162
rect 3110 3158 3114 3162
rect 3126 3158 3130 3162
rect 3174 3158 3178 3162
rect 3222 3158 3226 3162
rect 3278 3158 3282 3162
rect 3342 3158 3346 3162
rect 2710 3148 2714 3152
rect 2758 3148 2762 3152
rect 2918 3148 2922 3152
rect 2934 3148 2938 3152
rect 2998 3148 3002 3152
rect 3070 3148 3074 3152
rect 3134 3148 3138 3152
rect 3142 3148 3146 3152
rect 3190 3148 3194 3152
rect 3230 3148 3234 3152
rect 3262 3148 3266 3152
rect 3302 3148 3306 3152
rect 3318 3148 3322 3152
rect 3390 3158 3394 3162
rect 3438 3158 3442 3162
rect 3566 3158 3570 3162
rect 3590 3158 3594 3162
rect 3614 3158 3618 3162
rect 3702 3158 3706 3162
rect 3710 3158 3714 3162
rect 3358 3148 3362 3152
rect 3374 3148 3378 3152
rect 3446 3148 3450 3152
rect 3470 3148 3474 3152
rect 3558 3148 3562 3152
rect 3622 3148 3626 3152
rect 3654 3148 3658 3152
rect 3718 3148 3722 3152
rect 6 3138 10 3142
rect 70 3138 74 3142
rect 78 3138 82 3142
rect 214 3138 218 3142
rect 406 3138 410 3142
rect 582 3138 586 3142
rect 694 3138 698 3142
rect 710 3138 714 3142
rect 782 3138 786 3142
rect 822 3138 826 3142
rect 838 3138 842 3142
rect 902 3138 906 3142
rect 918 3138 922 3142
rect 942 3138 946 3142
rect 974 3138 978 3142
rect 1070 3138 1074 3142
rect 1126 3138 1130 3142
rect 1190 3138 1194 3142
rect 1262 3138 1266 3142
rect 1406 3138 1410 3142
rect 1470 3138 1474 3142
rect 1518 3138 1522 3142
rect 1526 3138 1530 3142
rect 1550 3138 1554 3142
rect 1686 3138 1690 3142
rect 1766 3138 1770 3142
rect 1774 3138 1778 3142
rect 1798 3138 1802 3142
rect 1822 3138 1826 3142
rect 1838 3138 1842 3142
rect 1886 3138 1890 3142
rect 1934 3138 1938 3142
rect 1942 3138 1946 3142
rect 1966 3138 1970 3142
rect 1990 3138 1994 3142
rect 2014 3138 2018 3142
rect 2046 3138 2050 3142
rect 2054 3138 2058 3142
rect 2110 3138 2114 3142
rect 2126 3138 2130 3142
rect 2134 3138 2138 3142
rect 2166 3138 2170 3142
rect 2222 3138 2226 3142
rect 2246 3138 2250 3142
rect 2254 3138 2258 3142
rect 2302 3138 2306 3142
rect 2310 3138 2314 3142
rect 2318 3138 2322 3142
rect 2326 3138 2330 3142
rect 2366 3138 2370 3142
rect 2398 3138 2402 3142
rect 2446 3138 2450 3142
rect 2454 3138 2458 3142
rect 2598 3138 2602 3142
rect 2630 3138 2634 3142
rect 2638 3138 2642 3142
rect 2686 3138 2690 3142
rect 2758 3138 2762 3142
rect 2934 3138 2938 3142
rect 2990 3138 2994 3142
rect 3014 3138 3018 3142
rect 3022 3138 3026 3142
rect 3078 3138 3082 3142
rect 3086 3138 3090 3142
rect 3150 3138 3154 3142
rect 3166 3138 3170 3142
rect 3206 3138 3210 3142
rect 3254 3138 3258 3142
rect 3326 3138 3330 3142
rect 3374 3138 3378 3142
rect 3398 3138 3402 3142
rect 3414 3138 3418 3142
rect 3438 3138 3442 3142
rect 3518 3138 3522 3142
rect 3574 3138 3578 3142
rect 3598 3138 3602 3142
rect 3662 3138 3666 3142
rect 3686 3138 3690 3142
rect 230 3128 234 3132
rect 422 3128 426 3132
rect 598 3128 602 3132
rect 934 3128 938 3132
rect 1086 3128 1090 3132
rect 1278 3128 1282 3132
rect 2350 3128 2354 3132
rect 2358 3128 2362 3132
rect 2470 3128 2474 3132
rect 2518 3128 2522 3132
rect 2566 3128 2570 3132
rect 2774 3128 2778 3132
rect 2862 3128 2866 3132
rect 3102 3128 3106 3132
rect 3166 3128 3170 3132
rect 3246 3128 3250 3132
rect 3286 3128 3290 3132
rect 3318 3128 3322 3132
rect 3390 3128 3394 3132
rect 3486 3128 3490 3132
rect 3502 3128 3506 3132
rect 3534 3128 3538 3132
rect 3646 3128 3650 3132
rect 3678 3128 3682 3132
rect 3742 3128 3746 3132
rect 3750 3128 3754 3132
rect 310 3118 314 3122
rect 502 3118 506 3122
rect 910 3118 914 3122
rect 1166 3118 1170 3122
rect 1182 3118 1186 3122
rect 1606 3118 1610 3122
rect 1630 3118 1634 3122
rect 1662 3118 1666 3122
rect 1790 3118 1794 3122
rect 2070 3118 2074 3122
rect 2118 3118 2122 3122
rect 2238 3118 2242 3122
rect 2462 3118 2466 3122
rect 2878 3118 2882 3122
rect 3046 3118 3050 3122
rect 3094 3118 3098 3122
rect 3158 3118 3162 3122
rect 3222 3118 3226 3122
rect 3238 3118 3242 3122
rect 3294 3118 3298 3122
rect 3310 3118 3314 3122
rect 3462 3118 3466 3122
rect 3478 3118 3482 3122
rect 3526 3118 3530 3122
rect 3558 3118 3562 3122
rect 3590 3118 3594 3122
rect 3638 3118 3642 3122
rect 3670 3118 3674 3122
rect 3702 3118 3706 3122
rect 850 3103 854 3107
rect 857 3103 861 3107
rect 1882 3103 1886 3107
rect 1889 3103 1893 3107
rect 2906 3103 2910 3107
rect 2913 3103 2917 3107
rect 766 3088 770 3092
rect 798 3088 802 3092
rect 822 3088 826 3092
rect 1094 3088 1098 3092
rect 1334 3088 1338 3092
rect 1518 3088 1522 3092
rect 1598 3088 1602 3092
rect 1622 3088 1626 3092
rect 1670 3088 1674 3092
rect 1718 3088 1722 3092
rect 1990 3088 1994 3092
rect 2054 3088 2058 3092
rect 2102 3088 2106 3092
rect 2190 3088 2194 3092
rect 2214 3088 2218 3092
rect 2310 3088 2314 3092
rect 2334 3088 2338 3092
rect 2350 3088 2354 3092
rect 2390 3088 2394 3092
rect 2478 3088 2482 3092
rect 2598 3088 2602 3092
rect 2630 3088 2634 3092
rect 2694 3088 2698 3092
rect 3094 3088 3098 3092
rect 3398 3088 3402 3092
rect 38 3078 42 3082
rect 118 3078 122 3082
rect 358 3078 362 3082
rect 582 3078 586 3082
rect 966 3078 970 3082
rect 1046 3078 1050 3082
rect 1246 3078 1250 3082
rect 1478 3078 1482 3082
rect 1870 3078 1874 3082
rect 1998 3078 2002 3082
rect 2014 3078 2018 3082
rect 2062 3078 2066 3082
rect 2206 3078 2210 3082
rect 2238 3078 2242 3082
rect 2302 3078 2306 3082
rect 2342 3078 2346 3082
rect 2382 3078 2386 3082
rect 2422 3078 2426 3082
rect 2806 3078 2810 3082
rect 3206 3078 3210 3082
rect 3214 3078 3218 3082
rect 3350 3078 3354 3082
rect 3486 3078 3490 3082
rect 3638 3078 3642 3082
rect 3710 3078 3714 3082
rect 3766 3078 3770 3082
rect 134 3068 138 3072
rect 206 3068 210 3072
rect 222 3068 226 3072
rect 230 3068 234 3072
rect 342 3068 346 3072
rect 439 3068 443 3072
rect 454 3068 458 3072
rect 566 3068 570 3072
rect 702 3068 706 3072
rect 742 3068 746 3072
rect 774 3068 778 3072
rect 862 3068 866 3072
rect 950 3068 954 3072
rect 1070 3068 1074 3072
rect 1086 3068 1090 3072
rect 1118 3068 1122 3072
rect 1134 3068 1138 3072
rect 1158 3068 1162 3072
rect 1262 3068 1266 3072
rect 1350 3068 1354 3072
rect 1438 3068 1442 3072
rect 1454 3068 1458 3072
rect 1486 3068 1490 3072
rect 1526 3068 1530 3072
rect 1574 3068 1578 3072
rect 1662 3068 1666 3072
rect 1694 3068 1698 3072
rect 1702 3068 1706 3072
rect 1718 3068 1722 3072
rect 1734 3068 1738 3072
rect 1758 3068 1762 3072
rect 1886 3068 1890 3072
rect 1974 3068 1978 3072
rect 2014 3068 2018 3072
rect 2046 3068 2050 3072
rect 2062 3068 2066 3072
rect 2086 3068 2090 3072
rect 22 3058 26 3062
rect 174 3058 178 3062
rect 222 3058 226 3062
rect 238 3058 242 3062
rect 294 3058 298 3062
rect 478 3058 482 3062
rect 486 3058 490 3062
rect 518 3058 522 3062
rect 622 3058 626 3062
rect 678 3058 682 3062
rect 694 3058 698 3062
rect 734 3058 738 3062
rect 750 3058 754 3062
rect 782 3058 786 3062
rect 806 3058 810 3062
rect 838 3058 842 3062
rect 854 3058 858 3062
rect 902 3058 906 3062
rect 1006 3058 1010 3062
rect 1078 3058 1082 3062
rect 1110 3058 1114 3062
rect 1206 3058 1210 3062
rect 1382 3058 1386 3062
rect 1414 3058 1418 3062
rect 1446 3058 1450 3062
rect 1462 3058 1466 3062
rect 1534 3058 1538 3062
rect 1550 3058 1554 3062
rect 1582 3058 1586 3062
rect 1614 3058 1618 3062
rect 1638 3058 1642 3062
rect 1694 3058 1698 3062
rect 1734 3058 1738 3062
rect 1830 3058 1834 3062
rect 1918 3058 1922 3062
rect 1998 3058 2002 3062
rect 2022 3058 2026 3062
rect 2038 3058 2042 3062
rect 2078 3058 2082 3062
rect 2118 3058 2122 3062
rect 2142 3068 2146 3072
rect 2134 3058 2138 3062
rect 2150 3058 2154 3062
rect 2166 3068 2170 3072
rect 2182 3068 2186 3072
rect 2222 3068 2226 3072
rect 2262 3068 2266 3072
rect 2294 3068 2298 3072
rect 2374 3068 2378 3072
rect 2470 3068 2474 3072
rect 2494 3068 2498 3072
rect 2502 3068 2506 3072
rect 2534 3068 2538 3072
rect 2582 3068 2586 3072
rect 2590 3068 2594 3072
rect 2622 3068 2626 3072
rect 2670 3068 2674 3072
rect 2678 3068 2682 3072
rect 2702 3068 2706 3072
rect 2822 3068 2826 3072
rect 2974 3068 2978 3072
rect 3054 3068 3058 3072
rect 3086 3068 3090 3072
rect 3118 3068 3122 3072
rect 3134 3068 3138 3072
rect 3214 3068 3218 3072
rect 3262 3068 3266 3072
rect 3270 3068 3274 3072
rect 3302 3068 3306 3072
rect 3374 3068 3378 3072
rect 3406 3068 3410 3072
rect 3454 3068 3458 3072
rect 3510 3068 3514 3072
rect 3638 3068 3642 3072
rect 3654 3068 3658 3072
rect 3670 3068 3674 3072
rect 3718 3068 3722 3072
rect 3734 3068 3738 3072
rect 2238 3058 2242 3062
rect 2254 3058 2258 3062
rect 2270 3058 2274 3062
rect 2286 3058 2290 3062
rect 2318 3058 2322 3062
rect 2366 3058 2370 3062
rect 2398 3058 2402 3062
rect 2430 3058 2434 3062
rect 2438 3058 2442 3062
rect 2462 3058 2466 3062
rect 2510 3058 2514 3062
rect 2614 3058 2618 3062
rect 2662 3058 2666 3062
rect 2702 3058 2706 3062
rect 2766 3058 2770 3062
rect 2870 3058 2874 3062
rect 3062 3058 3066 3062
rect 3078 3058 3082 3062
rect 3110 3058 3114 3062
rect 3182 3058 3186 3062
rect 3230 3058 3234 3062
rect 3254 3058 3258 3062
rect 3278 3058 3282 3062
rect 3294 3058 3298 3062
rect 3302 3058 3306 3062
rect 3334 3058 3338 3062
rect 3382 3058 3386 3062
rect 3430 3058 3434 3062
rect 3438 3058 3442 3062
rect 3462 3058 3466 3062
rect 3486 3058 3490 3062
rect 3502 3058 3506 3062
rect 3510 3058 3514 3062
rect 3558 3058 3562 3062
rect 3582 3058 3586 3062
rect 3622 3058 3626 3062
rect 3646 3058 3650 3062
rect 3662 3058 3666 3062
rect 3678 3058 3682 3062
rect 3694 3058 3698 3062
rect 3726 3058 3730 3062
rect 3750 3058 3754 3062
rect 182 3048 186 3052
rect 238 3048 242 3052
rect 254 3048 258 3052
rect 310 3050 314 3054
rect 534 3050 538 3054
rect 678 3048 682 3052
rect 766 3048 770 3052
rect 798 3048 802 3052
rect 838 3048 842 3052
rect 918 3050 922 3054
rect 1062 3048 1066 3052
rect 1094 3048 1098 3052
rect 1134 3048 1138 3052
rect 1294 3050 1298 3054
rect 1334 3048 1338 3052
rect 1350 3048 1354 3052
rect 1406 3048 1410 3052
rect 1430 3048 1434 3052
rect 1462 3048 1466 3052
rect 1502 3048 1506 3052
rect 1542 3048 1546 3052
rect 1598 3048 1602 3052
rect 1606 3048 1610 3052
rect 1670 3048 1674 3052
rect 1742 3048 1746 3052
rect 1758 3048 1762 3052
rect 1782 3048 1786 3052
rect 1934 3048 1938 3052
rect 1990 3048 1994 3052
rect 2094 3048 2098 3052
rect 2102 3048 2106 3052
rect 2134 3048 2138 3052
rect 2182 3048 2186 3052
rect 2198 3048 2202 3052
rect 2238 3048 2242 3052
rect 2270 3048 2274 3052
rect 2350 3048 2354 3052
rect 2446 3048 2450 3052
rect 2462 3048 2466 3052
rect 2478 3048 2482 3052
rect 2526 3048 2530 3052
rect 2566 3048 2570 3052
rect 2606 3048 2610 3052
rect 2646 3048 2650 3052
rect 2694 3048 2698 3052
rect 2854 3050 2858 3054
rect 3094 3048 3098 3052
rect 3142 3048 3146 3052
rect 3166 3048 3170 3052
rect 3238 3048 3242 3052
rect 3326 3048 3330 3052
rect 3366 3048 3370 3052
rect 3398 3048 3402 3052
rect 3446 3048 3450 3052
rect 3462 3048 3466 3052
rect 3478 3048 3482 3052
rect 3534 3048 3538 3052
rect 3566 3048 3570 3052
rect 3590 3048 3594 3052
rect 3742 3048 3746 3052
rect 6 3038 10 3042
rect 662 3038 666 3042
rect 1390 3038 1394 3042
rect 1422 3038 1426 3042
rect 1558 3038 1562 3042
rect 1622 3038 1626 3042
rect 2718 3038 2722 3042
rect 3126 3038 3130 3042
rect 3294 3038 3298 3042
rect 3518 3038 3522 3042
rect 3550 3038 3554 3042
rect 3582 3038 3586 3042
rect 310 3027 314 3031
rect 918 3027 922 3031
rect 1166 3028 1170 3032
rect 1294 3027 1298 3031
rect 1550 3028 1554 3032
rect 1766 3028 1770 3032
rect 2542 3028 2546 3032
rect 182 3018 186 3022
rect 494 3018 498 3022
rect 534 3018 538 3022
rect 1126 3018 1130 3022
rect 1382 3018 1386 3022
rect 1790 3018 1794 3022
rect 1934 3018 1938 3022
rect 2326 3018 2330 3022
rect 2726 3018 2730 3022
rect 2854 3018 2858 3022
rect 2918 3018 2922 3022
rect 3038 3018 3042 3022
rect 3062 3018 3066 3022
rect 3150 3018 3154 3022
rect 3254 3018 3258 3022
rect 3310 3018 3314 3022
rect 3558 3018 3562 3022
rect 3574 3018 3578 3022
rect 3622 3018 3626 3022
rect 3678 3018 3682 3022
rect 3758 3018 3762 3022
rect 346 3003 350 3007
rect 353 3003 357 3007
rect 1362 3003 1366 3007
rect 1369 3003 1373 3007
rect 2386 3003 2390 3007
rect 2393 3003 2397 3007
rect 3410 3003 3414 3007
rect 3417 3003 3421 3007
rect 86 2988 90 2992
rect 230 2988 234 2992
rect 526 2988 530 2992
rect 662 2988 666 2992
rect 686 2988 690 2992
rect 750 2988 754 2992
rect 782 2988 786 2992
rect 814 2988 818 2992
rect 918 2988 922 2992
rect 1006 2988 1010 2992
rect 1038 2988 1042 2992
rect 1446 2988 1450 2992
rect 1486 2988 1490 2992
rect 1574 2988 1578 2992
rect 1718 2988 1722 2992
rect 2126 2988 2130 2992
rect 2334 2988 2338 2992
rect 2414 2988 2418 2992
rect 2462 2988 2466 2992
rect 2726 2988 2730 2992
rect 3118 2988 3122 2992
rect 3462 2988 3466 2992
rect 366 2979 370 2983
rect 710 2978 714 2982
rect 1262 2978 1266 2982
rect 1870 2979 1874 2983
rect 2198 2978 2202 2982
rect 2902 2979 2906 2983
rect 2990 2979 2994 2983
rect 550 2968 554 2972
rect 654 2968 658 2972
rect 678 2968 682 2972
rect 742 2968 746 2972
rect 806 2968 810 2972
rect 894 2968 898 2972
rect 910 2968 914 2972
rect 966 2968 970 2972
rect 998 2968 1002 2972
rect 1230 2968 1234 2972
rect 1294 2968 1298 2972
rect 1318 2968 1322 2972
rect 1366 2968 1370 2972
rect 1494 2968 1498 2972
rect 1558 2968 1562 2972
rect 1582 2968 1586 2972
rect 1710 2968 1714 2972
rect 2094 2968 2098 2972
rect 3278 2968 3282 2972
rect 3334 2968 3338 2972
rect 3342 2968 3346 2972
rect 3454 2968 3458 2972
rect 3670 2968 3674 2972
rect 366 2956 370 2960
rect 510 2958 514 2962
rect 542 2958 546 2962
rect 566 2958 570 2962
rect 630 2958 634 2962
rect 638 2958 642 2962
rect 694 2958 698 2962
rect 758 2958 762 2962
rect 830 2958 834 2962
rect 934 2958 938 2962
rect 982 2958 986 2962
rect 1014 2958 1018 2962
rect 1038 2958 1042 2962
rect 1222 2958 1226 2962
rect 1278 2958 1282 2962
rect 1302 2958 1306 2962
rect 1382 2958 1386 2962
rect 1478 2958 1482 2962
rect 1526 2958 1530 2962
rect 1606 2958 1610 2962
rect 1622 2958 1626 2962
rect 1670 2958 1674 2962
rect 1678 2958 1682 2962
rect 1694 2958 1698 2962
rect 1726 2958 1730 2962
rect 22 2948 26 2952
rect 166 2948 170 2952
rect 342 2948 346 2952
rect 454 2948 458 2952
rect 526 2948 530 2952
rect 558 2948 562 2952
rect 598 2948 602 2952
rect 614 2948 618 2952
rect 646 2948 650 2952
rect 686 2948 690 2952
rect 726 2948 730 2952
rect 750 2948 754 2952
rect 766 2948 770 2952
rect 814 2948 818 2952
rect 846 2948 850 2952
rect 918 2948 922 2952
rect 950 2948 954 2952
rect 1006 2948 1010 2952
rect 1142 2948 1146 2952
rect 1206 2948 1210 2952
rect 1246 2948 1250 2952
rect 1286 2948 1290 2952
rect 1318 2948 1322 2952
rect 1406 2948 1410 2952
rect 1438 2948 1442 2952
rect 1470 2948 1474 2952
rect 1486 2948 1490 2952
rect 1534 2948 1538 2952
rect 1566 2948 1570 2952
rect 1590 2948 1594 2952
rect 1870 2956 1874 2960
rect 1974 2958 1978 2962
rect 2046 2958 2050 2962
rect 2054 2958 2058 2962
rect 2110 2958 2114 2962
rect 2142 2958 2146 2962
rect 2158 2958 2162 2962
rect 2214 2958 2218 2962
rect 2262 2958 2266 2962
rect 2430 2958 2434 2962
rect 2446 2958 2450 2962
rect 2478 2958 2482 2962
rect 1718 2948 1722 2952
rect 1782 2948 1786 2952
rect 1926 2948 1930 2952
rect 1982 2948 1986 2952
rect 2022 2948 2026 2952
rect 2030 2948 2034 2952
rect 2054 2948 2058 2952
rect 2070 2948 2074 2952
rect 2126 2948 2130 2952
rect 2158 2948 2162 2952
rect 2182 2948 2186 2952
rect 2222 2948 2226 2952
rect 2246 2948 2250 2952
rect 2270 2948 2274 2952
rect 2302 2948 2306 2952
rect 2310 2948 2314 2952
rect 2342 2948 2346 2952
rect 2350 2948 2354 2952
rect 2374 2948 2378 2952
rect 2430 2948 2434 2952
rect 2454 2948 2458 2952
rect 2478 2948 2482 2952
rect 2542 2958 2546 2962
rect 2726 2958 2730 2962
rect 2902 2956 2906 2960
rect 2926 2958 2930 2962
rect 2510 2948 2514 2952
rect 2558 2948 2562 2952
rect 2622 2948 2626 2952
rect 2710 2948 2714 2952
rect 2870 2948 2874 2952
rect 2990 2956 2994 2960
rect 3134 2958 3138 2962
rect 3158 2958 3162 2962
rect 3294 2958 3298 2962
rect 3318 2958 3322 2962
rect 3342 2958 3346 2962
rect 3350 2958 3354 2962
rect 3414 2958 3418 2962
rect 3502 2958 3506 2962
rect 3542 2958 3546 2962
rect 3654 2958 3658 2962
rect 3734 2958 3738 2962
rect 2974 2948 2978 2952
rect 3262 2948 3266 2952
rect 3286 2948 3290 2952
rect 3334 2948 3338 2952
rect 3382 2948 3386 2952
rect 3398 2948 3402 2952
rect 3446 2948 3450 2952
rect 3582 2948 3586 2952
rect 3614 2948 3618 2952
rect 3646 2948 3650 2952
rect 3662 2948 3666 2952
rect 3686 2948 3690 2952
rect 3726 2948 3730 2952
rect 3774 2948 3778 2952
rect 6 2938 10 2942
rect 30 2938 34 2942
rect 102 2938 106 2942
rect 174 2938 178 2942
rect 246 2938 250 2942
rect 310 2938 314 2942
rect 398 2938 402 2942
rect 534 2938 538 2942
rect 574 2938 578 2942
rect 606 2938 610 2942
rect 862 2938 866 2942
rect 870 2938 874 2942
rect 958 2938 962 2942
rect 982 2938 986 2942
rect 1086 2938 1090 2942
rect 1198 2938 1202 2942
rect 1214 2938 1218 2942
rect 1230 2938 1234 2942
rect 1310 2938 1314 2942
rect 1342 2938 1346 2942
rect 1398 2938 1402 2942
rect 1446 2938 1450 2942
rect 1462 2938 1466 2942
rect 1510 2938 1514 2942
rect 1542 2938 1546 2942
rect 1558 2938 1562 2942
rect 1630 2938 1634 2942
rect 1646 2938 1650 2942
rect 1654 2938 1658 2942
rect 1694 2938 1698 2942
rect 1838 2938 1842 2942
rect 1958 2938 1962 2942
rect 1990 2938 1994 2942
rect 2006 2938 2010 2942
rect 2014 2938 2018 2942
rect 2070 2938 2074 2942
rect 2134 2938 2138 2942
rect 2190 2938 2194 2942
rect 2238 2938 2242 2942
rect 2270 2938 2274 2942
rect 2294 2938 2298 2942
rect 2350 2938 2354 2942
rect 2382 2938 2386 2942
rect 2422 2938 2426 2942
rect 2454 2938 2458 2942
rect 2502 2938 2506 2942
rect 2534 2938 2538 2942
rect 2566 2938 2570 2942
rect 2581 2938 2585 2942
rect 2678 2938 2682 2942
rect 2750 2938 2754 2942
rect 2773 2938 2777 2942
rect 2870 2938 2874 2942
rect 3022 2938 3026 2942
rect 3150 2938 3154 2942
rect 3174 2938 3178 2942
rect 3182 2938 3186 2942
rect 3230 2938 3234 2942
rect 3254 2938 3258 2942
rect 3302 2938 3306 2942
rect 3318 2938 3322 2942
rect 3374 2938 3378 2942
rect 3390 2938 3394 2942
rect 3470 2938 3474 2942
rect 3518 2938 3522 2942
rect 3526 2938 3530 2942
rect 3542 2938 3546 2942
rect 3550 2938 3554 2942
rect 3558 2940 3562 2944
rect 3590 2938 3594 2942
rect 3630 2938 3634 2942
rect 3638 2938 3642 2942
rect 3734 2938 3738 2942
rect 414 2928 418 2932
rect 1102 2928 1106 2932
rect 1182 2928 1186 2932
rect 1422 2928 1426 2932
rect 1822 2928 1826 2932
rect 1998 2928 2002 2932
rect 2182 2928 2186 2932
rect 2222 2928 2226 2932
rect 2366 2928 2370 2932
rect 2398 2928 2402 2932
rect 2662 2928 2666 2932
rect 2766 2928 2770 2932
rect 2854 2928 2858 2932
rect 3038 2928 3042 2932
rect 3238 2928 3242 2932
rect 3358 2928 3362 2932
rect 3606 2928 3610 2932
rect 3702 2928 3706 2932
rect 3750 2928 3754 2932
rect 3758 2928 3762 2932
rect 86 2918 90 2922
rect 158 2918 162 2922
rect 494 2918 498 2922
rect 630 2918 634 2922
rect 886 2918 890 2922
rect 1366 2918 1370 2922
rect 1526 2918 1530 2922
rect 1638 2918 1642 2922
rect 1670 2918 1674 2922
rect 1742 2918 1746 2922
rect 1942 2918 1946 2922
rect 1974 2918 1978 2922
rect 2062 2918 2066 2922
rect 2254 2918 2258 2922
rect 2278 2918 2282 2922
rect 3142 2918 3146 2922
rect 3166 2918 3170 2922
rect 3214 2918 3218 2922
rect 3246 2918 3250 2922
rect 3278 2918 3282 2922
rect 3366 2918 3370 2922
rect 3574 2918 3578 2922
rect 3598 2918 3602 2922
rect 3662 2918 3666 2922
rect 3694 2918 3698 2922
rect 3710 2918 3714 2922
rect 3766 2918 3770 2922
rect 850 2903 854 2907
rect 857 2903 861 2907
rect 1882 2903 1886 2907
rect 1889 2903 1893 2907
rect 2906 2903 2910 2907
rect 2913 2903 2917 2907
rect 630 2888 634 2892
rect 662 2888 666 2892
rect 750 2888 754 2892
rect 806 2888 810 2892
rect 878 2888 882 2892
rect 934 2888 938 2892
rect 982 2888 986 2892
rect 1462 2888 1466 2892
rect 1710 2888 1714 2892
rect 1966 2888 1970 2892
rect 2046 2888 2050 2892
rect 2118 2888 2122 2892
rect 2342 2888 2346 2892
rect 2462 2888 2466 2892
rect 2486 2888 2490 2892
rect 2614 2888 2618 2892
rect 2662 2888 2666 2892
rect 2758 2888 2762 2892
rect 2798 2888 2802 2892
rect 3270 2888 3274 2892
rect 3454 2888 3458 2892
rect 3566 2888 3570 2892
rect 30 2878 34 2882
rect 94 2878 98 2882
rect 334 2878 338 2882
rect 526 2878 530 2882
rect 606 2878 610 2882
rect 622 2878 626 2882
rect 742 2878 746 2882
rect 1182 2878 1186 2882
rect 1350 2878 1354 2882
rect 1406 2878 1410 2882
rect 1422 2878 1426 2882
rect 1606 2878 1610 2882
rect 1742 2878 1746 2882
rect 1854 2878 1858 2882
rect 2094 2878 2098 2882
rect 2126 2878 2130 2882
rect 2302 2878 2306 2882
rect 2422 2878 2426 2882
rect 2542 2878 2546 2882
rect 2622 2878 2626 2882
rect 2694 2878 2698 2882
rect 2742 2878 2746 2882
rect 54 2868 58 2872
rect 118 2868 122 2872
rect 214 2868 218 2872
rect 222 2868 226 2872
rect 238 2868 242 2872
rect 318 2868 322 2872
rect 374 2868 378 2872
rect 510 2868 514 2872
rect 670 2868 674 2872
rect 742 2868 746 2872
rect 766 2868 770 2872
rect 774 2868 778 2872
rect 830 2868 834 2872
rect 862 2868 866 2872
rect 910 2868 914 2872
rect 998 2868 1002 2872
rect 1014 2868 1018 2872
rect 1030 2868 1034 2872
rect 1094 2868 1098 2872
rect 1166 2868 1170 2872
rect 1263 2868 1267 2872
rect 1294 2868 1298 2872
rect 1310 2868 1314 2872
rect 1350 2868 1354 2872
rect 1366 2868 1370 2872
rect 1414 2868 1418 2872
rect 1422 2868 1426 2872
rect 1438 2868 1442 2872
rect 1446 2868 1450 2872
rect 1494 2868 1498 2872
rect 1510 2868 1514 2872
rect 1622 2868 1626 2872
rect 1702 2868 1706 2872
rect 1718 2868 1722 2872
rect 1870 2868 1874 2872
rect 2014 2868 2018 2872
rect 2022 2868 2026 2872
rect 2070 2868 2074 2872
rect 2110 2868 2114 2872
rect 2126 2868 2130 2872
rect 2150 2868 2154 2872
rect 2190 2868 2194 2872
rect 2222 2868 2226 2872
rect 2286 2868 2290 2872
rect 2294 2868 2298 2872
rect 2318 2868 2322 2872
rect 2334 2868 2338 2872
rect 2366 2868 2370 2872
rect 2398 2868 2402 2872
rect 2406 2868 2410 2872
rect 2478 2868 2482 2872
rect 2558 2868 2562 2872
rect 22 2858 26 2862
rect 46 2858 50 2862
rect 62 2858 66 2862
rect 110 2858 114 2862
rect 126 2858 130 2862
rect 222 2858 226 2862
rect 270 2858 274 2862
rect 462 2858 466 2862
rect 646 2858 650 2862
rect 678 2858 682 2862
rect 694 2858 698 2862
rect 718 2858 722 2862
rect 782 2858 786 2862
rect 822 2858 826 2862
rect 854 2858 858 2862
rect 902 2858 906 2862
rect 918 2858 922 2862
rect 974 2858 978 2862
rect 1022 2858 1026 2862
rect 1054 2858 1058 2862
rect 1070 2858 1074 2862
rect 1086 2858 1090 2862
rect 1126 2858 1130 2862
rect 1222 2858 1226 2862
rect 1334 2858 1338 2862
rect 1382 2858 1386 2862
rect 1470 2858 1474 2862
rect 1654 2858 1658 2862
rect 1662 2858 1666 2862
rect 1694 2858 1698 2862
rect 1734 2858 1738 2862
rect 1758 2858 1762 2862
rect 1918 2858 1922 2862
rect 1926 2858 1930 2862
rect 1982 2858 1986 2862
rect 2062 2858 2066 2862
rect 2078 2858 2082 2862
rect 2102 2858 2106 2862
rect 2142 2858 2146 2862
rect 2166 2858 2170 2862
rect 2214 2858 2218 2862
rect 2230 2858 2234 2862
rect 2254 2858 2258 2862
rect 2278 2858 2282 2862
rect 2326 2858 2330 2862
rect 2390 2858 2394 2862
rect 2438 2858 2442 2862
rect 2446 2858 2450 2862
rect 2518 2858 2522 2862
rect 2566 2858 2570 2862
rect 2582 2868 2586 2872
rect 2606 2868 2610 2872
rect 2622 2868 2626 2872
rect 2646 2868 2650 2872
rect 2686 2868 2690 2872
rect 2718 2868 2722 2872
rect 2806 2878 2810 2882
rect 2822 2878 2826 2882
rect 2902 2878 2906 2882
rect 2990 2878 2994 2882
rect 3262 2878 3266 2882
rect 3318 2878 3322 2882
rect 3374 2878 3378 2882
rect 3422 2878 3426 2882
rect 3654 2878 3658 2882
rect 3726 2878 3730 2882
rect 3766 2878 3770 2882
rect 2766 2868 2770 2872
rect 2774 2868 2778 2872
rect 2918 2868 2922 2872
rect 3118 2868 3122 2872
rect 3150 2868 3154 2872
rect 3198 2868 3202 2872
rect 3206 2868 3210 2872
rect 3254 2868 3258 2872
rect 3278 2868 3282 2872
rect 3310 2868 3314 2872
rect 3382 2868 3386 2872
rect 3470 2868 3474 2872
rect 3518 2868 3522 2872
rect 3526 2868 3530 2872
rect 3582 2868 3586 2872
rect 3614 2868 3618 2872
rect 3638 2868 3642 2872
rect 3654 2868 3658 2872
rect 3686 2868 3690 2872
rect 3718 2868 3722 2872
rect 2590 2858 2594 2862
rect 2598 2858 2602 2862
rect 2638 2858 2642 2862
rect 2678 2858 2682 2862
rect 2710 2858 2714 2862
rect 2726 2858 2730 2862
rect 2774 2858 2778 2862
rect 2966 2858 2970 2862
rect 3030 2858 3034 2862
rect 3062 2858 3066 2862
rect 3094 2858 3098 2862
rect 3126 2858 3130 2862
rect 3150 2858 3154 2862
rect 3334 2858 3338 2862
rect 3358 2858 3362 2862
rect 3390 2858 3394 2862
rect 3550 2858 3554 2862
rect 3590 2858 3594 2862
rect 3670 2858 3674 2862
rect 3742 2858 3746 2862
rect 62 2848 66 2852
rect 78 2848 82 2852
rect 126 2848 130 2852
rect 142 2848 146 2852
rect 246 2848 250 2852
rect 286 2850 290 2854
rect 478 2850 482 2854
rect 662 2848 666 2852
rect 726 2848 730 2852
rect 750 2848 754 2852
rect 798 2848 802 2852
rect 806 2848 810 2852
rect 838 2848 842 2852
rect 886 2848 890 2852
rect 982 2848 986 2852
rect 1006 2848 1010 2852
rect 1054 2848 1058 2852
rect 1134 2850 1138 2854
rect 1270 2848 1274 2852
rect 1294 2848 1298 2852
rect 1342 2848 1346 2852
rect 1398 2848 1402 2852
rect 1454 2848 1458 2852
rect 1670 2848 1674 2852
rect 1902 2850 1906 2854
rect 2038 2848 2042 2852
rect 2158 2848 2162 2852
rect 2166 2848 2170 2852
rect 2198 2848 2202 2852
rect 2262 2848 2266 2852
rect 2310 2848 2314 2852
rect 2342 2848 2346 2852
rect 2374 2848 2378 2852
rect 2502 2848 2506 2852
rect 2550 2848 2554 2852
rect 2654 2848 2658 2852
rect 2662 2848 2666 2852
rect 2694 2848 2698 2852
rect 2950 2850 2954 2854
rect 3022 2848 3026 2852
rect 3054 2848 3058 2852
rect 3086 2848 3090 2852
rect 3142 2848 3146 2852
rect 3294 2848 3298 2852
rect 3326 2848 3330 2852
rect 3406 2848 3410 2852
rect 3462 2848 3466 2852
rect 3542 2848 3546 2852
rect 3606 2848 3610 2852
rect 3694 2848 3698 2852
rect 6 2838 10 2842
rect 430 2838 434 2842
rect 710 2838 714 2842
rect 782 2838 786 2842
rect 1046 2838 1050 2842
rect 1342 2838 1346 2842
rect 1470 2838 1474 2842
rect 2998 2838 3002 2842
rect 3038 2838 3042 2842
rect 3070 2838 3074 2842
rect 3102 2838 3106 2842
rect 3342 2838 3346 2842
rect 3446 2838 3450 2842
rect 3590 2838 3594 2842
rect 286 2827 290 2831
rect 478 2827 482 2831
rect 1334 2828 1338 2832
rect 1902 2827 1906 2831
rect 3238 2828 3242 2832
rect 3366 2828 3370 2832
rect 94 2818 98 2822
rect 158 2818 162 2822
rect 854 2818 858 2822
rect 958 2818 962 2822
rect 1134 2818 1138 2822
rect 1302 2818 1306 2822
rect 1486 2818 1490 2822
rect 1502 2818 1506 2822
rect 1526 2818 1530 2822
rect 1670 2818 1674 2822
rect 1774 2818 1778 2822
rect 2006 2818 2010 2822
rect 2278 2818 2282 2822
rect 2534 2818 2538 2822
rect 2790 2818 2794 2822
rect 2950 2818 2954 2822
rect 3046 2818 3050 2822
rect 3078 2818 3082 2822
rect 3094 2818 3098 2822
rect 3126 2818 3130 2822
rect 3350 2818 3354 2822
rect 3390 2818 3394 2822
rect 3502 2818 3506 2822
rect 3534 2818 3538 2822
rect 3750 2818 3754 2822
rect 346 2803 350 2807
rect 353 2803 357 2807
rect 1362 2803 1366 2807
rect 1369 2803 1373 2807
rect 2386 2803 2390 2807
rect 2393 2803 2397 2807
rect 3410 2803 3414 2807
rect 3417 2803 3421 2807
rect 182 2788 186 2792
rect 358 2788 362 2792
rect 414 2788 418 2792
rect 590 2788 594 2792
rect 678 2788 682 2792
rect 742 2788 746 2792
rect 774 2788 778 2792
rect 982 2788 986 2792
rect 1046 2788 1050 2792
rect 1110 2788 1114 2792
rect 1134 2788 1138 2792
rect 1278 2788 1282 2792
rect 1414 2788 1418 2792
rect 1454 2788 1458 2792
rect 1518 2788 1522 2792
rect 1662 2788 1666 2792
rect 1846 2788 1850 2792
rect 2078 2788 2082 2792
rect 2222 2788 2226 2792
rect 2302 2788 2306 2792
rect 2422 2788 2426 2792
rect 2462 2788 2466 2792
rect 2814 2788 2818 2792
rect 2926 2788 2930 2792
rect 3070 2788 3074 2792
rect 3254 2788 3258 2792
rect 646 2778 650 2782
rect 606 2768 610 2772
rect 806 2778 810 2782
rect 926 2778 930 2782
rect 2590 2779 2594 2783
rect 3126 2779 3130 2783
rect 3438 2778 3442 2782
rect 718 2768 722 2772
rect 782 2768 786 2772
rect 798 2768 802 2772
rect 942 2768 946 2772
rect 1422 2768 1426 2772
rect 1710 2768 1714 2772
rect 1734 2768 1738 2772
rect 1990 2768 1994 2772
rect 3710 2768 3714 2772
rect 3726 2768 3730 2772
rect 182 2758 186 2762
rect 358 2758 362 2762
rect 414 2758 418 2762
rect 614 2758 618 2762
rect 662 2758 666 2762
rect 702 2758 706 2762
rect 758 2758 762 2762
rect 766 2758 770 2762
rect 798 2758 802 2762
rect 838 2758 842 2762
rect 862 2758 866 2762
rect 878 2758 882 2762
rect 910 2758 914 2762
rect 998 2758 1002 2762
rect 1278 2758 1282 2762
rect 1334 2758 1338 2762
rect 1406 2758 1410 2762
rect 1662 2758 1666 2762
rect 1758 2758 1762 2762
rect 1782 2758 1786 2762
rect 1822 2758 1826 2762
rect 174 2748 178 2752
rect 342 2748 346 2752
rect 422 2748 426 2752
rect 606 2748 610 2752
rect 622 2748 626 2752
rect 678 2748 682 2752
rect 710 2748 714 2752
rect 742 2748 746 2752
rect 774 2748 778 2752
rect 806 2748 810 2752
rect 838 2748 842 2752
rect 894 2748 898 2752
rect 926 2748 930 2752
rect 942 2748 946 2752
rect 990 2748 994 2752
rect 998 2748 1002 2752
rect 1014 2748 1018 2752
rect 1030 2748 1034 2752
rect 1062 2748 1066 2752
rect 1094 2748 1098 2752
rect 1230 2748 1234 2752
rect 1326 2748 1330 2752
rect 1366 2748 1370 2752
rect 1422 2748 1426 2752
rect 1438 2748 1442 2752
rect 1470 2748 1474 2752
rect 1510 2748 1514 2752
rect 1558 2748 1562 2752
rect 1654 2748 1658 2752
rect 1686 2748 1690 2752
rect 1718 2748 1722 2752
rect 1726 2748 1730 2752
rect 1742 2748 1746 2752
rect 1910 2758 1914 2762
rect 2006 2758 2010 2762
rect 2222 2758 2226 2762
rect 2262 2758 2266 2762
rect 2310 2758 2314 2762
rect 2342 2758 2346 2762
rect 2374 2758 2378 2762
rect 2590 2756 2594 2760
rect 2630 2758 2634 2762
rect 2734 2758 2738 2762
rect 2774 2758 2778 2762
rect 2790 2758 2794 2762
rect 2830 2758 2834 2762
rect 3070 2758 3074 2762
rect 3078 2758 3082 2762
rect 1846 2748 1850 2752
rect 1910 2748 1914 2752
rect 1934 2748 1938 2752
rect 1942 2748 1946 2752
rect 1990 2748 1994 2752
rect 2030 2748 2034 2752
rect 2062 2748 2066 2752
rect 2214 2748 2218 2752
rect 2262 2748 2266 2752
rect 2286 2748 2290 2752
rect 2318 2748 2322 2752
rect 2358 2748 2362 2752
rect 2414 2748 2418 2752
rect 2454 2748 2458 2752
rect 2606 2748 2610 2752
rect 2646 2748 2650 2752
rect 2662 2748 2666 2752
rect 2718 2748 2722 2752
rect 2742 2748 2746 2752
rect 2790 2748 2794 2752
rect 2798 2748 2802 2752
rect 2846 2748 2850 2752
rect 2862 2748 2866 2752
rect 2870 2748 2874 2752
rect 2910 2748 2914 2752
rect 2966 2748 2970 2752
rect 3126 2756 3130 2760
rect 3294 2758 3298 2762
rect 3470 2758 3474 2762
rect 3542 2758 3546 2762
rect 3598 2758 3602 2762
rect 3694 2758 3698 2762
rect 3758 2758 3762 2762
rect 3110 2748 3114 2752
rect 3262 2748 3266 2752
rect 3270 2748 3274 2752
rect 3358 2748 3362 2752
rect 3382 2748 3386 2752
rect 3454 2748 3458 2752
rect 3502 2748 3506 2752
rect 3558 2748 3562 2752
rect 3566 2748 3570 2752
rect 3614 2748 3618 2752
rect 3630 2748 3634 2752
rect 3670 2748 3674 2752
rect 3702 2748 3706 2752
rect 6 2738 10 2742
rect 134 2738 138 2742
rect 310 2738 314 2742
rect 462 2738 466 2742
rect 559 2738 563 2742
rect 574 2738 578 2742
rect 638 2738 642 2742
rect 670 2738 674 2742
rect 734 2738 738 2742
rect 830 2738 834 2742
rect 902 2738 906 2742
rect 934 2738 938 2742
rect 958 2738 962 2742
rect 990 2738 994 2742
rect 1022 2738 1026 2742
rect 1230 2738 1234 2742
rect 1318 2738 1322 2742
rect 1350 2738 1354 2742
rect 1398 2738 1402 2742
rect 1478 2738 1482 2742
rect 1494 2738 1498 2742
rect 1614 2738 1618 2742
rect 1694 2738 1698 2742
rect 1710 2738 1714 2742
rect 1774 2738 1778 2742
rect 1798 2738 1802 2742
rect 1806 2738 1810 2742
rect 1878 2738 1882 2742
rect 1894 2738 1898 2742
rect 2014 2738 2018 2742
rect 2038 2738 2042 2742
rect 2046 2738 2050 2742
rect 2070 2738 2074 2742
rect 2174 2738 2178 2742
rect 2254 2738 2258 2742
rect 2286 2738 2290 2742
rect 2294 2738 2298 2742
rect 2334 2738 2338 2742
rect 2366 2738 2370 2742
rect 2382 2738 2386 2742
rect 2398 2738 2402 2742
rect 2438 2738 2442 2742
rect 2558 2738 2562 2742
rect 2638 2738 2642 2742
rect 2654 2738 2658 2742
rect 2670 2738 2674 2742
rect 2694 2738 2698 2742
rect 2798 2738 2802 2742
rect 2806 2738 2810 2742
rect 2854 2738 2858 2742
rect 2870 2738 2874 2742
rect 3022 2738 3026 2742
rect 3158 2738 3162 2742
rect 3270 2738 3274 2742
rect 3302 2738 3306 2742
rect 3390 2738 3394 2742
rect 3430 2738 3434 2742
rect 3446 2738 3450 2742
rect 3494 2738 3498 2742
rect 3518 2738 3522 2742
rect 3566 2738 3570 2742
rect 3622 2738 3626 2742
rect 3662 2738 3666 2742
rect 3742 2738 3746 2742
rect 3758 2738 3762 2742
rect 3774 2738 3778 2742
rect 118 2728 122 2732
rect 294 2728 298 2732
rect 478 2728 482 2732
rect 966 2728 970 2732
rect 1214 2728 1218 2732
rect 1302 2728 1306 2732
rect 1598 2728 1602 2732
rect 1862 2728 1866 2732
rect 1958 2728 1962 2732
rect 2158 2728 2162 2732
rect 2422 2728 2426 2732
rect 2542 2728 2546 2732
rect 2686 2728 2690 2732
rect 2766 2728 2770 2732
rect 2838 2728 2842 2732
rect 2894 2728 2898 2732
rect 3006 2728 3010 2732
rect 3174 2728 3178 2732
rect 3374 2728 3378 2732
rect 3406 2728 3410 2732
rect 3534 2728 3538 2732
rect 3590 2728 3594 2732
rect 3750 2728 3754 2732
rect 214 2718 218 2722
rect 582 2718 586 2722
rect 630 2718 634 2722
rect 878 2718 882 2722
rect 1046 2718 1050 2722
rect 1078 2718 1082 2722
rect 1310 2718 1314 2722
rect 1342 2718 1346 2722
rect 1486 2718 1490 2722
rect 1790 2718 1794 2722
rect 2022 2718 2026 2722
rect 2246 2718 2250 2722
rect 2678 2718 2682 2722
rect 2702 2718 2706 2722
rect 2758 2718 2762 2722
rect 2926 2718 2930 2722
rect 3294 2718 3298 2722
rect 3334 2718 3338 2722
rect 3398 2718 3402 2722
rect 3486 2718 3490 2722
rect 3526 2718 3530 2722
rect 3542 2718 3546 2722
rect 3582 2718 3586 2722
rect 3598 2718 3602 2722
rect 3686 2718 3690 2722
rect 850 2703 854 2707
rect 857 2703 861 2707
rect 1882 2703 1886 2707
rect 1889 2703 1893 2707
rect 2906 2703 2910 2707
rect 2913 2703 2917 2707
rect 374 2688 378 2692
rect 478 2688 482 2692
rect 518 2688 522 2692
rect 694 2688 698 2692
rect 750 2688 754 2692
rect 830 2688 834 2692
rect 854 2688 858 2692
rect 966 2688 970 2692
rect 1054 2688 1058 2692
rect 1110 2688 1114 2692
rect 1142 2688 1146 2692
rect 1486 2688 1490 2692
rect 1638 2688 1642 2692
rect 1718 2688 1722 2692
rect 1782 2688 1786 2692
rect 1854 2688 1858 2692
rect 2110 2688 2114 2692
rect 2134 2688 2138 2692
rect 2206 2688 2210 2692
rect 2438 2688 2442 2692
rect 2462 2688 2466 2692
rect 2638 2688 2642 2692
rect 2734 2688 2738 2692
rect 2822 2688 2826 2692
rect 230 2678 234 2682
rect 366 2678 370 2682
rect 582 2678 586 2682
rect 662 2678 666 2682
rect 758 2678 762 2682
rect 974 2678 978 2682
rect 1030 2678 1034 2682
rect 1046 2678 1050 2682
rect 1086 2678 1090 2682
rect 1222 2678 1226 2682
rect 1406 2678 1410 2682
rect 1526 2678 1530 2682
rect 1534 2678 1538 2682
rect 1566 2678 1570 2682
rect 1726 2678 1730 2682
rect 1758 2678 1762 2682
rect 1998 2678 2002 2682
rect 2094 2678 2098 2682
rect 2102 2678 2106 2682
rect 2214 2678 2218 2682
rect 2446 2678 2450 2682
rect 2542 2678 2546 2682
rect 2646 2678 2650 2682
rect 2702 2678 2706 2682
rect 2902 2678 2906 2682
rect 2926 2678 2930 2682
rect 3046 2678 3050 2682
rect 3174 2678 3178 2682
rect 3238 2678 3242 2682
rect 3286 2678 3290 2682
rect 3326 2678 3330 2682
rect 3350 2678 3354 2682
rect 3406 2678 3410 2682
rect 3462 2678 3466 2682
rect 3486 2678 3490 2682
rect 3590 2678 3594 2682
rect 3630 2678 3634 2682
rect 3670 2678 3674 2682
rect 3702 2678 3706 2682
rect 3710 2678 3714 2682
rect 78 2668 82 2672
rect 214 2668 218 2672
rect 318 2668 322 2672
rect 342 2668 346 2672
rect 398 2668 402 2672
rect 430 2668 434 2672
rect 438 2668 442 2672
rect 454 2668 458 2672
rect 542 2668 546 2672
rect 614 2668 618 2672
rect 630 2668 634 2672
rect 646 2668 650 2672
rect 670 2668 674 2672
rect 702 2668 706 2672
rect 742 2668 746 2672
rect 766 2668 770 2672
rect 782 2668 786 2672
rect 798 2668 802 2672
rect 806 2668 810 2672
rect 838 2668 842 2672
rect 862 2668 866 2672
rect 918 2668 922 2672
rect 950 2668 954 2672
rect 982 2668 986 2672
rect 998 2668 1002 2672
rect 1014 2668 1018 2672
rect 1078 2668 1082 2672
rect 1126 2668 1130 2672
rect 1238 2668 1242 2672
rect 1390 2668 1394 2672
rect 1574 2668 1578 2672
rect 1590 2668 1594 2672
rect 1622 2668 1626 2672
rect 1662 2668 1666 2672
rect 1678 2668 1682 2672
rect 1694 2668 1698 2672
rect 1710 2668 1714 2672
rect 1734 2668 1738 2672
rect 1750 2668 1754 2672
rect 1774 2668 1778 2672
rect 1806 2668 1810 2672
rect 1814 2668 1818 2672
rect 1838 2668 1842 2672
rect 1902 2668 1906 2672
rect 2014 2668 2018 2672
rect 2118 2668 2122 2672
rect 2142 2668 2146 2672
rect 2174 2668 2178 2672
rect 2198 2668 2202 2672
rect 2222 2668 2226 2672
rect 2238 2668 2242 2672
rect 2254 2668 2258 2672
rect 2310 2668 2314 2672
rect 2342 2668 2346 2672
rect 2382 2668 2386 2672
rect 2390 2668 2394 2672
rect 2558 2668 2562 2672
rect 2630 2668 2634 2672
rect 2686 2668 2690 2672
rect 2742 2668 2746 2672
rect 2782 2668 2786 2672
rect 2790 2668 2794 2672
rect 2846 2668 2850 2672
rect 2862 2668 2866 2672
rect 2878 2668 2882 2672
rect 2950 2668 2954 2672
rect 3030 2668 3034 2672
rect 3166 2668 3170 2672
rect 3190 2668 3194 2672
rect 3230 2668 3234 2672
rect 3262 2668 3266 2672
rect 3270 2668 3274 2672
rect 3294 2668 3298 2672
rect 3470 2668 3474 2672
rect 3486 2668 3490 2672
rect 3614 2668 3618 2672
rect 3638 2668 3642 2672
rect 6 2658 10 2662
rect 174 2658 178 2662
rect 311 2658 315 2662
rect 350 2658 354 2662
rect 390 2658 394 2662
rect 406 2658 410 2662
rect 422 2658 426 2662
rect 462 2658 466 2662
rect 502 2658 506 2662
rect 534 2658 538 2662
rect 566 2658 570 2662
rect 598 2658 602 2662
rect 622 2658 626 2662
rect 638 2658 642 2662
rect 678 2658 682 2662
rect 710 2658 714 2662
rect 726 2658 730 2662
rect 742 2658 746 2662
rect 774 2658 778 2662
rect 790 2658 794 2662
rect 814 2658 818 2662
rect 830 2658 834 2662
rect 902 2658 906 2662
rect 926 2658 930 2662
rect 942 2658 946 2662
rect 958 2658 962 2662
rect 990 2658 994 2662
rect 1006 2658 1010 2662
rect 1030 2658 1034 2662
rect 1038 2658 1042 2662
rect 1070 2658 1074 2662
rect 1102 2658 1106 2662
rect 1286 2658 1290 2662
rect 182 2650 186 2654
rect 374 2648 378 2652
rect 406 2648 410 2652
rect 478 2648 482 2652
rect 486 2648 490 2652
rect 510 2648 514 2652
rect 574 2648 578 2652
rect 582 2648 586 2652
rect 694 2648 698 2652
rect 726 2648 730 2652
rect 910 2648 914 2652
rect 942 2648 946 2652
rect 1054 2648 1058 2652
rect 1270 2650 1274 2654
rect 1446 2658 1450 2662
rect 1550 2658 1554 2662
rect 1582 2658 1586 2662
rect 1614 2658 1618 2662
rect 1654 2658 1658 2662
rect 1686 2658 1690 2662
rect 1702 2658 1706 2662
rect 1798 2658 1802 2662
rect 1822 2658 1826 2662
rect 1878 2658 1882 2662
rect 1958 2658 1962 2662
rect 2094 2658 2098 2662
rect 2118 2658 2122 2662
rect 2150 2658 2154 2662
rect 2190 2658 2194 2662
rect 2230 2658 2234 2662
rect 2262 2658 2266 2662
rect 2366 2658 2370 2662
rect 2374 2658 2378 2662
rect 2422 2658 2426 2662
rect 2430 2658 2434 2662
rect 2606 2658 2610 2662
rect 2662 2658 2666 2662
rect 2694 2658 2698 2662
rect 2718 2658 2722 2662
rect 2758 2658 2762 2662
rect 2774 2658 2778 2662
rect 2798 2658 2802 2662
rect 2814 2658 2818 2662
rect 2838 2658 2842 2662
rect 2854 2658 2858 2662
rect 2886 2658 2890 2662
rect 2902 2658 2906 2662
rect 2942 2658 2946 2662
rect 3086 2658 3090 2662
rect 3158 2658 3162 2662
rect 3198 2658 3202 2662
rect 3222 2658 3226 2662
rect 3254 2658 3258 2662
rect 3326 2658 3330 2662
rect 3350 2658 3354 2662
rect 3366 2658 3370 2662
rect 3382 2658 3386 2662
rect 3422 2658 3426 2662
rect 3446 2658 3450 2662
rect 3470 2658 3474 2662
rect 3542 2658 3546 2662
rect 3566 2658 3570 2662
rect 3574 2658 3578 2662
rect 3606 2658 3610 2662
rect 3630 2658 3634 2662
rect 3662 2658 3666 2662
rect 3702 2658 3706 2662
rect 3734 2658 3738 2662
rect 1334 2648 1338 2652
rect 1358 2650 1362 2654
rect 1510 2648 1514 2652
rect 1630 2648 1634 2652
rect 1638 2648 1642 2652
rect 1670 2648 1674 2652
rect 1782 2648 1786 2652
rect 1830 2648 1834 2652
rect 1862 2648 1866 2652
rect 2062 2648 2066 2652
rect 2166 2648 2170 2652
rect 2246 2648 2250 2652
rect 2278 2648 2282 2652
rect 2318 2648 2322 2652
rect 2350 2648 2354 2652
rect 2422 2648 2426 2652
rect 2590 2650 2594 2654
rect 2758 2648 2762 2652
rect 2814 2648 2818 2652
rect 2822 2648 2826 2652
rect 2958 2648 2962 2652
rect 2998 2650 3002 2654
rect 3142 2648 3146 2652
rect 3206 2648 3210 2652
rect 3398 2648 3402 2652
rect 3518 2648 3522 2652
rect 3558 2648 3562 2652
rect 3590 2648 3594 2652
rect 3630 2648 3634 2652
rect 3662 2648 3666 2652
rect 3774 2648 3778 2652
rect 494 2638 498 2642
rect 558 2638 562 2642
rect 846 2638 850 2642
rect 894 2638 898 2642
rect 2774 2638 2778 2642
rect 3126 2638 3130 2642
rect 3342 2638 3346 2642
rect 3534 2638 3538 2642
rect 182 2627 186 2631
rect 446 2628 450 2632
rect 1270 2627 1274 2631
rect 2302 2628 2306 2632
rect 2590 2627 2594 2631
rect 2670 2628 2674 2632
rect 3566 2628 3570 2632
rect 62 2618 66 2622
rect 134 2618 138 2622
rect 566 2618 570 2622
rect 886 2618 890 2622
rect 1358 2618 1362 2622
rect 1518 2618 1522 2622
rect 1598 2618 1602 2622
rect 1766 2618 1770 2622
rect 1918 2618 1922 2622
rect 2062 2618 2066 2622
rect 2150 2618 2154 2622
rect 2182 2618 2186 2622
rect 2998 2618 3002 2622
rect 3158 2618 3162 2622
rect 3174 2618 3178 2622
rect 3222 2618 3226 2622
rect 3254 2618 3258 2622
rect 3286 2618 3290 2622
rect 3382 2618 3386 2622
rect 3438 2618 3442 2622
rect 3502 2618 3506 2622
rect 3526 2618 3530 2622
rect 3678 2618 3682 2622
rect 3734 2618 3738 2622
rect 346 2603 350 2607
rect 353 2603 357 2607
rect 1362 2603 1366 2607
rect 1369 2603 1373 2607
rect 2386 2603 2390 2607
rect 2393 2603 2397 2607
rect 3410 2603 3414 2607
rect 3417 2603 3421 2607
rect 182 2588 186 2592
rect 358 2588 362 2592
rect 614 2588 618 2592
rect 758 2588 762 2592
rect 822 2588 826 2592
rect 902 2588 906 2592
rect 974 2588 978 2592
rect 1046 2588 1050 2592
rect 1086 2588 1090 2592
rect 1222 2588 1226 2592
rect 1550 2588 1554 2592
rect 1582 2588 1586 2592
rect 1806 2588 1810 2592
rect 1942 2588 1946 2592
rect 2166 2588 2170 2592
rect 2310 2588 2314 2592
rect 2422 2588 2426 2592
rect 2534 2588 2538 2592
rect 2742 2588 2746 2592
rect 2806 2588 2810 2592
rect 2878 2588 2882 2592
rect 2934 2588 2938 2592
rect 2990 2588 2994 2592
rect 3710 2588 3714 2592
rect 534 2579 538 2583
rect 694 2578 698 2582
rect 934 2578 938 2582
rect 1350 2579 1354 2583
rect 2070 2579 2074 2583
rect 2382 2578 2386 2582
rect 2582 2578 2586 2582
rect 6 2568 10 2572
rect 702 2568 706 2572
rect 766 2568 770 2572
rect 830 2568 834 2572
rect 1542 2568 1546 2572
rect 1790 2568 1794 2572
rect 1814 2568 1818 2572
rect 2718 2568 2722 2572
rect 3182 2568 3186 2572
rect 182 2558 186 2562
rect 358 2558 362 2562
rect 534 2556 538 2560
rect 574 2558 578 2562
rect 646 2558 650 2562
rect 654 2558 658 2562
rect 686 2558 690 2562
rect 718 2558 722 2562
rect 750 2558 754 2562
rect 790 2558 794 2562
rect 806 2558 810 2562
rect 814 2558 818 2562
rect 886 2558 890 2562
rect 1006 2558 1010 2562
rect 1118 2558 1122 2562
rect 1166 2558 1170 2562
rect 1278 2558 1282 2562
rect 1350 2556 1354 2560
rect 1510 2558 1514 2562
rect 1526 2558 1530 2562
rect 1558 2558 1562 2562
rect 1582 2558 1586 2562
rect 1830 2558 1834 2562
rect 1886 2558 1890 2562
rect 2070 2556 2074 2560
rect 2110 2558 2114 2562
rect 2142 2558 2146 2562
rect 2310 2558 2314 2562
rect 2358 2558 2362 2562
rect 2366 2558 2370 2562
rect 2438 2558 2442 2562
rect 2446 2558 2450 2562
rect 2478 2558 2482 2562
rect 2550 2558 2554 2562
rect 2566 2558 2570 2562
rect 2598 2558 2602 2562
rect 2606 2558 2610 2562
rect 2646 2558 2650 2562
rect 2662 2558 2666 2562
rect 2670 2558 2674 2562
rect 2702 2558 2706 2562
rect 2822 2558 2826 2562
rect 2854 2558 2858 2562
rect 2862 2558 2866 2562
rect 174 2548 178 2552
rect 182 2548 186 2552
rect 254 2548 258 2552
rect 358 2548 362 2552
rect 446 2548 450 2552
rect 574 2548 578 2552
rect 630 2548 634 2552
rect 670 2548 674 2552
rect 702 2548 706 2552
rect 734 2548 738 2552
rect 758 2548 762 2552
rect 790 2548 794 2552
rect 822 2548 826 2552
rect 870 2548 874 2552
rect 886 2548 890 2552
rect 918 2548 922 2552
rect 958 2548 962 2552
rect 990 2548 994 2552
rect 1054 2548 1058 2552
rect 1078 2548 1082 2552
rect 1134 2548 1138 2552
rect 1150 2548 1154 2552
rect 1182 2548 1186 2552
rect 1206 2548 1210 2552
rect 1222 2548 1226 2552
rect 1246 2548 1250 2552
rect 1262 2548 1266 2552
rect 1382 2548 1386 2552
rect 1510 2548 1514 2552
rect 1550 2548 1554 2552
rect 1582 2548 1586 2552
rect 1758 2548 1762 2552
rect 1766 2548 1770 2552
rect 1798 2548 1802 2552
rect 1822 2548 1826 2552
rect 1862 2548 1866 2552
rect 1910 2548 1914 2552
rect 1982 2548 1986 2552
rect 2094 2548 2098 2552
rect 2134 2548 2138 2552
rect 2206 2548 2210 2552
rect 2342 2548 2346 2552
rect 2382 2548 2386 2552
rect 2422 2548 2426 2552
rect 2454 2548 2458 2552
rect 2502 2548 2506 2552
rect 2510 2548 2514 2552
rect 2542 2548 2546 2552
rect 2574 2548 2578 2552
rect 2638 2548 2642 2552
rect 2646 2548 2650 2552
rect 2670 2548 2674 2552
rect 2686 2548 2690 2552
rect 2718 2548 2722 2552
rect 2742 2548 2746 2552
rect 2790 2548 2794 2552
rect 2806 2548 2810 2552
rect 2830 2548 2834 2552
rect 2862 2548 2866 2552
rect 2878 2548 2882 2552
rect 2910 2548 2914 2552
rect 2958 2558 2962 2562
rect 3030 2558 3034 2562
rect 3086 2558 3090 2562
rect 3110 2558 3114 2562
rect 3214 2558 3218 2562
rect 3254 2558 3258 2562
rect 3318 2558 3322 2562
rect 3398 2558 3402 2562
rect 3494 2558 3498 2562
rect 3518 2558 3522 2562
rect 3542 2558 3546 2562
rect 3590 2558 3594 2562
rect 3614 2558 3618 2562
rect 3646 2558 3650 2562
rect 3694 2558 3698 2562
rect 3742 2558 3746 2562
rect 3758 2558 3762 2562
rect 3774 2558 3778 2562
rect 2974 2548 2978 2552
rect 3006 2548 3010 2552
rect 3038 2548 3042 2552
rect 134 2538 138 2542
rect 310 2538 314 2542
rect 502 2538 506 2542
rect 598 2538 602 2542
rect 606 2538 610 2542
rect 622 2538 626 2542
rect 638 2538 642 2542
rect 678 2538 682 2542
rect 718 2538 722 2542
rect 742 2538 746 2542
rect 782 2538 786 2542
rect 862 2538 866 2542
rect 1054 2538 1058 2542
rect 1062 2538 1066 2542
rect 1102 2538 1106 2542
rect 1126 2538 1130 2542
rect 1158 2538 1162 2542
rect 1190 2538 1194 2542
rect 1198 2538 1202 2542
rect 1230 2538 1234 2542
rect 1238 2538 1242 2542
rect 1254 2538 1258 2542
rect 1270 2538 1274 2542
rect 1294 2538 1298 2542
rect 1382 2538 1386 2542
rect 1494 2538 1498 2542
rect 3118 2548 3122 2552
rect 3158 2548 3162 2552
rect 3174 2548 3178 2552
rect 3294 2548 3298 2552
rect 3342 2548 3346 2552
rect 3366 2548 3370 2552
rect 3374 2548 3378 2552
rect 3446 2548 3450 2552
rect 3478 2548 3482 2552
rect 3574 2548 3578 2552
rect 3614 2548 3618 2552
rect 3638 2548 3642 2552
rect 3670 2548 3674 2552
rect 3686 2548 3690 2552
rect 3726 2548 3730 2552
rect 3758 2548 3762 2552
rect 1630 2538 1634 2542
rect 1774 2538 1778 2542
rect 1798 2538 1802 2542
rect 1910 2538 1914 2542
rect 1918 2538 1922 2542
rect 2038 2538 2042 2542
rect 2126 2538 2130 2542
rect 2262 2538 2266 2542
rect 2334 2538 2338 2542
rect 2350 2538 2354 2542
rect 2390 2538 2394 2542
rect 2406 2538 2410 2542
rect 2470 2538 2474 2542
rect 2502 2538 2506 2542
rect 2518 2538 2522 2542
rect 2542 2538 2546 2542
rect 2574 2538 2578 2542
rect 2630 2538 2634 2542
rect 2638 2538 2642 2542
rect 2694 2538 2698 2542
rect 2726 2538 2730 2542
rect 2734 2538 2738 2542
rect 2782 2538 2786 2542
rect 2798 2538 2802 2542
rect 2830 2538 2834 2542
rect 2886 2538 2890 2542
rect 2894 2538 2898 2542
rect 2926 2538 2930 2542
rect 2982 2538 2986 2542
rect 2998 2538 3002 2542
rect 3046 2538 3050 2542
rect 3062 2538 3066 2542
rect 3070 2538 3074 2542
rect 3094 2538 3098 2542
rect 3174 2538 3178 2542
rect 3198 2538 3202 2542
rect 3230 2538 3234 2542
rect 3238 2538 3242 2542
rect 3262 2538 3266 2542
rect 3286 2538 3290 2542
rect 3294 2538 3298 2542
rect 3502 2538 3506 2542
rect 3526 2538 3530 2542
rect 3542 2538 3546 2542
rect 3622 2538 3626 2542
rect 3638 2538 3642 2542
rect 3662 2538 3666 2542
rect 3670 2538 3674 2542
rect 3718 2538 3722 2542
rect 3734 2538 3738 2542
rect 3750 2538 3754 2542
rect 118 2528 122 2532
rect 294 2528 298 2532
rect 406 2528 410 2532
rect 486 2528 490 2532
rect 1094 2528 1098 2532
rect 1398 2528 1402 2532
rect 1646 2528 1650 2532
rect 1734 2528 1738 2532
rect 1758 2528 1762 2532
rect 1838 2528 1842 2532
rect 1846 2528 1850 2532
rect 2022 2528 2026 2532
rect 2150 2528 2154 2532
rect 2246 2528 2250 2532
rect 2534 2528 2538 2532
rect 2766 2528 2770 2532
rect 3062 2528 3066 2532
rect 3158 2528 3162 2532
rect 3286 2528 3290 2532
rect 3326 2528 3330 2532
rect 3342 2528 3346 2532
rect 3406 2528 3410 2532
rect 3462 2528 3466 2532
rect 3702 2528 3706 2532
rect 214 2518 218 2522
rect 654 2518 658 2522
rect 1070 2518 1074 2522
rect 1118 2518 1122 2522
rect 1150 2518 1154 2522
rect 1166 2518 1170 2522
rect 1286 2518 1290 2522
rect 1502 2518 1506 2522
rect 1926 2518 1930 2522
rect 2118 2518 2122 2522
rect 2606 2518 2610 2522
rect 2902 2518 2906 2522
rect 3030 2518 3034 2522
rect 3086 2518 3090 2522
rect 3142 2518 3146 2522
rect 3318 2518 3322 2522
rect 3334 2518 3338 2522
rect 3398 2518 3402 2522
rect 3414 2518 3418 2522
rect 3494 2518 3498 2522
rect 3518 2518 3522 2522
rect 3542 2518 3546 2522
rect 3654 2518 3658 2522
rect 850 2503 854 2507
rect 857 2503 861 2507
rect 1882 2503 1886 2507
rect 1889 2503 1893 2507
rect 2906 2503 2910 2507
rect 2913 2503 2917 2507
rect 462 2488 466 2492
rect 710 2488 714 2492
rect 942 2488 946 2492
rect 974 2488 978 2492
rect 1062 2488 1066 2492
rect 1222 2488 1226 2492
rect 1230 2488 1234 2492
rect 1342 2488 1346 2492
rect 1398 2488 1402 2492
rect 1542 2488 1546 2492
rect 1558 2488 1562 2492
rect 1638 2488 1642 2492
rect 1766 2488 1770 2492
rect 1878 2488 1882 2492
rect 2014 2488 2018 2492
rect 2054 2488 2058 2492
rect 2182 2488 2186 2492
rect 2230 2488 2234 2492
rect 2262 2488 2266 2492
rect 2278 2488 2282 2492
rect 2334 2488 2338 2492
rect 2382 2488 2386 2492
rect 2534 2488 2538 2492
rect 2750 2488 2754 2492
rect 2798 2488 2802 2492
rect 2854 2488 2858 2492
rect 2934 2488 2938 2492
rect 3134 2488 3138 2492
rect 3166 2488 3170 2492
rect 3190 2488 3194 2492
rect 3222 2488 3226 2492
rect 3278 2488 3282 2492
rect 3630 2488 3634 2492
rect 6 2478 10 2482
rect 174 2478 178 2482
rect 366 2478 370 2482
rect 550 2478 554 2482
rect 998 2478 1002 2482
rect 1094 2478 1098 2482
rect 1102 2478 1106 2482
rect 1118 2478 1122 2482
rect 1150 2478 1154 2482
rect 1182 2478 1186 2482
rect 1254 2478 1258 2482
rect 1726 2478 1730 2482
rect 1734 2478 1738 2482
rect 1750 2478 1754 2482
rect 1758 2478 1762 2482
rect 1790 2478 1794 2482
rect 2062 2478 2066 2482
rect 2206 2478 2210 2482
rect 2222 2478 2226 2482
rect 2286 2478 2290 2482
rect 2310 2478 2314 2482
rect 2342 2478 2346 2482
rect 2350 2478 2354 2482
rect 2374 2478 2378 2482
rect 2422 2478 2426 2482
rect 2486 2478 2490 2482
rect 2614 2478 2618 2482
rect 2806 2478 2810 2482
rect 2838 2478 2842 2482
rect 2846 2478 2850 2482
rect 2926 2478 2930 2482
rect 2982 2478 2986 2482
rect 3014 2478 3018 2482
rect 3094 2478 3098 2482
rect 3142 2478 3146 2482
rect 3198 2478 3202 2482
rect 3230 2478 3234 2482
rect 3238 2478 3242 2482
rect 3286 2478 3290 2482
rect 3294 2478 3298 2482
rect 3310 2478 3314 2482
rect 3398 2478 3402 2482
rect 3566 2478 3570 2482
rect 3590 2478 3594 2482
rect 30 2468 34 2472
rect 54 2468 58 2472
rect 93 2468 97 2472
rect 190 2468 194 2472
rect 382 2468 386 2472
rect 454 2468 458 2472
rect 534 2468 538 2472
rect 631 2468 635 2472
rect 718 2468 722 2472
rect 806 2468 810 2472
rect 838 2468 842 2472
rect 894 2468 898 2472
rect 926 2468 930 2472
rect 934 2468 938 2472
rect 966 2468 970 2472
rect 990 2468 994 2472
rect 1014 2468 1018 2472
rect 1038 2468 1042 2472
rect 1086 2468 1090 2472
rect 1110 2468 1114 2472
rect 1142 2468 1146 2472
rect 1166 2468 1170 2472
rect 1206 2468 1210 2472
rect 1270 2468 1274 2472
rect 1286 2468 1290 2472
rect 1406 2468 1410 2472
rect 1446 2468 1450 2472
rect 1518 2468 1522 2472
rect 1550 2468 1554 2472
rect 1574 2468 1578 2472
rect 1582 2468 1586 2472
rect 1654 2468 1658 2472
rect 1686 2468 1690 2472
rect 1718 2468 1722 2472
rect 1774 2468 1778 2472
rect 1846 2468 1850 2472
rect 1854 2468 1858 2472
rect 1894 2468 1898 2472
rect 1950 2468 1954 2472
rect 1958 2468 1962 2472
rect 2006 2468 2010 2472
rect 2038 2468 2042 2472
rect 2070 2468 2074 2472
rect 2102 2468 2106 2472
rect 2150 2468 2154 2472
rect 2158 2468 2162 2472
rect 2310 2468 2314 2472
rect 2390 2468 2394 2472
rect 2430 2468 2434 2472
rect 2446 2468 2450 2472
rect 2494 2468 2498 2472
rect 2510 2468 2514 2472
rect 2630 2468 2634 2472
rect 2710 2468 2714 2472
rect 2726 2468 2730 2472
rect 2734 2468 2738 2472
rect 2758 2468 2762 2472
rect 2790 2468 2794 2472
rect 2814 2468 2818 2472
rect 2862 2468 2866 2472
rect 2886 2468 2890 2472
rect 2902 2468 2906 2472
rect 2942 2468 2946 2472
rect 2958 2468 2962 2472
rect 2998 2468 3002 2472
rect 3014 2468 3018 2472
rect 3062 2468 3066 2472
rect 3070 2468 3074 2472
rect 3126 2468 3130 2472
rect 3150 2468 3154 2472
rect 3182 2468 3186 2472
rect 3214 2468 3218 2472
rect 3238 2468 3242 2472
rect 3262 2468 3266 2472
rect 3366 2468 3370 2472
rect 3390 2468 3394 2472
rect 3398 2468 3402 2472
rect 3414 2468 3418 2472
rect 3646 2468 3650 2472
rect 3694 2468 3698 2472
rect 3702 2468 3706 2472
rect 3750 2468 3754 2472
rect 22 2458 26 2462
rect 46 2458 50 2462
rect 54 2458 58 2462
rect 238 2458 242 2462
rect 382 2458 386 2462
rect 430 2458 434 2462
rect 494 2458 498 2462
rect 654 2458 658 2462
rect 678 2458 682 2462
rect 686 2458 690 2462
rect 694 2458 698 2462
rect 734 2458 738 2462
rect 750 2458 754 2462
rect 774 2458 778 2462
rect 790 2458 794 2462
rect 814 2458 818 2462
rect 830 2458 834 2462
rect 886 2458 890 2462
rect 902 2458 906 2462
rect 918 2458 922 2462
rect 942 2458 946 2462
rect 958 2458 962 2462
rect 1014 2458 1018 2462
rect 1038 2458 1042 2462
rect 1070 2458 1074 2462
rect 1118 2458 1122 2462
rect 1134 2458 1138 2462
rect 1142 2458 1146 2462
rect 1174 2458 1178 2462
rect 1198 2458 1202 2462
rect 1278 2458 1282 2462
rect 1438 2458 1442 2462
rect 1526 2458 1530 2462
rect 1542 2458 1546 2462
rect 1662 2458 1666 2462
rect 1670 2458 1674 2462
rect 1694 2458 1698 2462
rect 1710 2458 1714 2462
rect 1814 2458 1818 2462
rect 1846 2458 1850 2462
rect 1854 2458 1858 2462
rect 1942 2458 1946 2462
rect 1966 2458 1970 2462
rect 2030 2458 2034 2462
rect 2046 2458 2050 2462
rect 2078 2458 2082 2462
rect 2126 2458 2130 2462
rect 2166 2458 2170 2462
rect 2190 2458 2194 2462
rect 2238 2458 2242 2462
rect 2246 2458 2250 2462
rect 2318 2458 2322 2462
rect 2366 2458 2370 2462
rect 2454 2458 2458 2462
rect 2502 2458 2506 2462
rect 2574 2458 2578 2462
rect 2670 2458 2674 2462
rect 2718 2458 2722 2462
rect 2782 2458 2786 2462
rect 2814 2458 2818 2462
rect 2870 2458 2874 2462
rect 2894 2458 2898 2462
rect 2950 2458 2954 2462
rect 2966 2458 2970 2462
rect 2990 2458 2994 2462
rect 3030 2458 3034 2462
rect 3110 2458 3114 2462
rect 3118 2458 3122 2462
rect 3174 2458 3178 2462
rect 3206 2458 3210 2462
rect 3254 2458 3258 2462
rect 3302 2458 3306 2462
rect 3326 2458 3330 2462
rect 3342 2458 3346 2462
rect 3350 2458 3354 2462
rect 3374 2458 3378 2462
rect 3414 2458 3418 2462
rect 3446 2458 3450 2462
rect 3486 2458 3490 2462
rect 3518 2458 3522 2462
rect 3550 2458 3554 2462
rect 3582 2458 3586 2462
rect 3606 2458 3610 2462
rect 3614 2458 3618 2462
rect 62 2448 66 2452
rect 78 2448 82 2452
rect 222 2450 226 2454
rect 286 2448 290 2452
rect 414 2450 418 2454
rect 486 2448 490 2452
rect 646 2448 650 2452
rect 782 2448 786 2452
rect 814 2448 818 2452
rect 974 2448 978 2452
rect 1222 2448 1226 2452
rect 1230 2448 1234 2452
rect 1558 2448 1562 2452
rect 1678 2448 1682 2452
rect 1822 2448 1826 2452
rect 1926 2448 1930 2452
rect 1982 2448 1986 2452
rect 2078 2448 2082 2452
rect 2118 2448 2122 2452
rect 2182 2448 2186 2452
rect 2470 2448 2474 2452
rect 2662 2450 2666 2454
rect 2702 2448 2706 2452
rect 2758 2448 2762 2452
rect 2774 2448 2778 2452
rect 2878 2448 2882 2452
rect 2982 2448 2986 2452
rect 3022 2448 3026 2452
rect 3086 2448 3090 2452
rect 3166 2448 3170 2452
rect 3278 2448 3282 2452
rect 3358 2448 3362 2452
rect 3390 2448 3394 2452
rect 3462 2448 3466 2452
rect 3494 2448 3498 2452
rect 3526 2448 3530 2452
rect 3550 2448 3554 2452
rect 638 2438 642 2442
rect 766 2438 770 2442
rect 790 2438 794 2442
rect 870 2438 874 2442
rect 1206 2438 1210 2442
rect 1422 2438 1426 2442
rect 1694 2438 1698 2442
rect 2366 2438 2370 2442
rect 3038 2438 3042 2442
rect 3478 2438 3482 2442
rect 3510 2438 3514 2442
rect 3542 2438 3546 2442
rect 918 2428 922 2432
rect 2662 2427 2666 2431
rect 3054 2428 3058 2432
rect 3446 2428 3450 2432
rect 222 2418 226 2422
rect 414 2418 418 2422
rect 486 2418 490 2422
rect 630 2418 634 2422
rect 654 2418 658 2422
rect 1502 2418 1506 2422
rect 1638 2418 1642 2422
rect 2518 2418 2522 2422
rect 2838 2418 2842 2422
rect 3030 2418 3034 2422
rect 3078 2418 3082 2422
rect 3110 2418 3114 2422
rect 3470 2418 3474 2422
rect 3518 2418 3522 2422
rect 3550 2418 3554 2422
rect 3582 2418 3586 2422
rect 3606 2418 3610 2422
rect 3670 2418 3674 2422
rect 3734 2418 3738 2422
rect 346 2403 350 2407
rect 353 2403 357 2407
rect 1362 2403 1366 2407
rect 1369 2403 1373 2407
rect 2386 2403 2390 2407
rect 2393 2403 2397 2407
rect 3410 2403 3414 2407
rect 3417 2403 3421 2407
rect 206 2388 210 2392
rect 246 2388 250 2392
rect 470 2388 474 2392
rect 494 2388 498 2392
rect 558 2388 562 2392
rect 638 2388 642 2392
rect 838 2388 842 2392
rect 982 2388 986 2392
rect 1006 2388 1010 2392
rect 1062 2388 1066 2392
rect 1254 2388 1258 2392
rect 1326 2388 1330 2392
rect 1726 2388 1730 2392
rect 1742 2388 1746 2392
rect 1758 2388 1762 2392
rect 1990 2388 1994 2392
rect 2046 2388 2050 2392
rect 2222 2388 2226 2392
rect 2262 2388 2266 2392
rect 2294 2388 2298 2392
rect 2750 2388 2754 2392
rect 2814 2388 2818 2392
rect 3046 2388 3050 2392
rect 3622 2388 3626 2392
rect 446 2378 450 2382
rect 606 2378 610 2382
rect 30 2368 34 2372
rect 526 2368 530 2372
rect 614 2368 618 2372
rect 686 2368 690 2372
rect 1190 2379 1194 2383
rect 1510 2379 1514 2383
rect 2390 2379 2394 2383
rect 758 2368 762 2372
rect 2078 2368 2082 2372
rect 3438 2368 3442 2372
rect 3670 2378 3674 2382
rect 3614 2368 3618 2372
rect 3702 2368 3706 2372
rect 3742 2368 3746 2372
rect 206 2358 210 2362
rect 246 2358 250 2362
rect 510 2358 514 2362
rect 542 2358 546 2362
rect 590 2358 594 2362
rect 598 2358 602 2362
rect 670 2358 674 2362
rect 702 2358 706 2362
rect 742 2358 746 2362
rect 790 2358 794 2362
rect 822 2358 826 2362
rect 950 2358 954 2362
rect 1030 2358 1034 2362
rect 1190 2356 1194 2360
rect 1510 2356 1514 2360
rect 1558 2358 1562 2362
rect 1574 2358 1578 2362
rect 1606 2358 1610 2362
rect 22 2348 26 2352
rect 206 2348 210 2352
rect 238 2348 242 2352
rect 350 2348 354 2352
rect 454 2348 458 2352
rect 486 2348 490 2352
rect 526 2348 530 2352
rect 606 2348 610 2352
rect 654 2348 658 2352
rect 686 2348 690 2352
rect 718 2348 722 2352
rect 750 2348 754 2352
rect 798 2348 802 2352
rect 822 2348 826 2352
rect 894 2348 898 2352
rect 910 2348 914 2352
rect 926 2348 930 2352
rect 966 2348 970 2352
rect 990 2348 994 2352
rect 1030 2348 1034 2352
rect 1198 2348 1202 2352
rect 1270 2348 1274 2352
rect 1294 2348 1298 2352
rect 1310 2348 1314 2352
rect 1334 2348 1338 2352
rect 1422 2348 1426 2352
rect 1558 2348 1562 2352
rect 1590 2348 1594 2352
rect 1670 2358 1674 2362
rect 1798 2358 1802 2362
rect 1822 2358 1826 2362
rect 1926 2358 1930 2362
rect 2030 2358 2034 2362
rect 2062 2358 2066 2362
rect 2222 2358 2226 2362
rect 2310 2358 2314 2362
rect 2390 2356 2394 2360
rect 2534 2358 2538 2362
rect 2662 2358 2666 2362
rect 3046 2358 3050 2362
rect 3150 2358 3154 2362
rect 3230 2358 3234 2362
rect 3406 2358 3410 2362
rect 3454 2358 3458 2362
rect 3462 2358 3466 2362
rect 3542 2358 3546 2362
rect 3598 2358 3602 2362
rect 3630 2358 3634 2362
rect 3686 2358 3690 2362
rect 3718 2358 3722 2362
rect 3750 2358 3754 2362
rect 1654 2348 1658 2352
rect 1670 2348 1674 2352
rect 1694 2348 1698 2352
rect 1782 2348 1786 2352
rect 1790 2348 1794 2352
rect 1830 2348 1834 2352
rect 1838 2348 1842 2352
rect 1854 2348 1858 2352
rect 1870 2348 1874 2352
rect 1886 2348 1890 2352
rect 1918 2348 1922 2352
rect 1942 2348 1946 2352
rect 2014 2348 2018 2352
rect 2030 2348 2034 2352
rect 2038 2348 2042 2352
rect 2222 2348 2226 2352
rect 2246 2348 2250 2352
rect 2278 2348 2282 2352
rect 2326 2348 2330 2352
rect 2366 2348 2370 2352
rect 2478 2348 2482 2352
rect 2550 2348 2554 2352
rect 2582 2348 2586 2352
rect 2646 2348 2650 2352
rect 2662 2348 2666 2352
rect 2678 2348 2682 2352
rect 2686 2348 2690 2352
rect 2702 2348 2706 2352
rect 2718 2348 2722 2352
rect 2734 2348 2738 2352
rect 2750 2348 2754 2352
rect 2798 2348 2802 2352
rect 2838 2348 2842 2352
rect 2870 2348 2874 2352
rect 3030 2348 3034 2352
rect 3070 2348 3074 2352
rect 3118 2348 3122 2352
rect 3174 2348 3178 2352
rect 3206 2348 3210 2352
rect 3262 2348 3266 2352
rect 3294 2348 3298 2352
rect 3326 2348 3330 2352
rect 3342 2348 3346 2352
rect 3350 2348 3354 2352
rect 3374 2348 3378 2352
rect 3390 2348 3394 2352
rect 3446 2348 3450 2352
rect 3470 2348 3474 2352
rect 3510 2348 3514 2352
rect 3526 2348 3530 2352
rect 3566 2348 3570 2352
rect 3582 2348 3586 2352
rect 3614 2348 3618 2352
rect 3654 2348 3658 2352
rect 3670 2348 3674 2352
rect 3710 2348 3714 2352
rect 3742 2348 3746 2352
rect 6 2338 10 2342
rect 158 2338 162 2342
rect 294 2338 298 2342
rect 438 2338 442 2342
rect 486 2338 490 2342
rect 518 2338 522 2342
rect 550 2338 554 2342
rect 566 2338 570 2342
rect 582 2338 586 2342
rect 662 2338 666 2342
rect 678 2338 682 2342
rect 710 2338 714 2342
rect 774 2338 778 2342
rect 790 2338 794 2342
rect 798 2338 802 2342
rect 862 2338 866 2342
rect 886 2338 890 2342
rect 902 2338 906 2342
rect 918 2338 922 2342
rect 1046 2338 1050 2342
rect 1158 2338 1162 2342
rect 1246 2338 1250 2342
rect 1278 2338 1282 2342
rect 1286 2338 1290 2342
rect 1302 2338 1306 2342
rect 1318 2338 1322 2342
rect 1478 2338 1482 2342
rect 1550 2338 1554 2342
rect 1582 2338 1586 2342
rect 1630 2338 1634 2342
rect 1662 2338 1666 2342
rect 1686 2338 1690 2342
rect 1718 2338 1722 2342
rect 1774 2338 1778 2342
rect 1806 2338 1810 2342
rect 1846 2338 1850 2342
rect 1950 2338 1954 2342
rect 1974 2338 1978 2342
rect 2006 2338 2010 2342
rect 2038 2338 2042 2342
rect 2174 2338 2178 2342
rect 2318 2338 2322 2342
rect 2334 2338 2338 2342
rect 2422 2338 2426 2342
rect 2542 2338 2546 2342
rect 2558 2338 2562 2342
rect 2606 2338 2610 2342
rect 2638 2338 2642 2342
rect 2654 2338 2658 2342
rect 2694 2338 2698 2342
rect 2734 2338 2738 2342
rect 2790 2338 2794 2342
rect 2806 2338 2810 2342
rect 2846 2338 2850 2342
rect 2862 2338 2866 2342
rect 2870 2338 2874 2342
rect 2998 2338 3002 2342
rect 3078 2338 3082 2342
rect 3126 2338 3130 2342
rect 3134 2338 3138 2342
rect 3174 2338 3178 2342
rect 3182 2338 3186 2342
rect 3198 2338 3202 2342
rect 3206 2338 3210 2342
rect 3230 2338 3234 2342
rect 3254 2338 3258 2342
rect 3262 2338 3266 2342
rect 3286 2338 3290 2342
rect 3598 2338 3602 2342
rect 3702 2338 3706 2342
rect 142 2328 146 2332
rect 310 2328 314 2332
rect 430 2328 434 2332
rect 934 2328 938 2332
rect 974 2328 978 2332
rect 1142 2328 1146 2332
rect 1230 2328 1234 2332
rect 1334 2328 1338 2332
rect 1374 2328 1378 2332
rect 1382 2328 1386 2332
rect 1462 2328 1466 2332
rect 1734 2328 1738 2332
rect 1750 2328 1754 2332
rect 1766 2328 1770 2332
rect 1814 2328 1818 2332
rect 1854 2328 1858 2332
rect 1870 2328 1874 2332
rect 1982 2328 1986 2332
rect 1998 2328 2002 2332
rect 2158 2328 2162 2332
rect 2438 2328 2442 2332
rect 2566 2328 2570 2332
rect 2622 2328 2626 2332
rect 2718 2328 2722 2332
rect 2774 2328 2778 2332
rect 2822 2328 2826 2332
rect 2982 2328 2986 2332
rect 3094 2328 3098 2332
rect 3158 2328 3162 2332
rect 3198 2328 3202 2332
rect 3238 2328 3242 2332
rect 3270 2328 3274 2332
rect 3334 2328 3338 2332
rect 3358 2328 3362 2332
rect 3494 2328 3498 2332
rect 3550 2328 3554 2332
rect 3638 2328 3642 2332
rect 390 2318 394 2322
rect 734 2318 738 2322
rect 838 2318 842 2322
rect 1038 2318 1042 2322
rect 1638 2318 1642 2322
rect 2518 2318 2522 2322
rect 2598 2318 2602 2322
rect 3102 2318 3106 2322
rect 3150 2318 3154 2322
rect 3230 2318 3234 2322
rect 3414 2318 3418 2322
rect 3486 2318 3490 2322
rect 3542 2318 3546 2322
rect 3734 2318 3738 2322
rect 850 2303 854 2307
rect 857 2303 861 2307
rect 1882 2303 1886 2307
rect 1889 2303 1893 2307
rect 2906 2303 2910 2307
rect 2913 2303 2917 2307
rect 486 2288 490 2292
rect 662 2288 666 2292
rect 926 2288 930 2292
rect 1022 2288 1026 2292
rect 1102 2288 1106 2292
rect 1166 2288 1170 2292
rect 1190 2288 1194 2292
rect 1222 2288 1226 2292
rect 1462 2288 1466 2292
rect 1518 2288 1522 2292
rect 1702 2288 1706 2292
rect 1846 2288 1850 2292
rect 1934 2288 1938 2292
rect 1982 2288 1986 2292
rect 2382 2288 2386 2292
rect 2590 2288 2594 2292
rect 2862 2288 2866 2292
rect 2894 2288 2898 2292
rect 2950 2288 2954 2292
rect 3006 2288 3010 2292
rect 3222 2288 3226 2292
rect 3566 2288 3570 2292
rect 326 2278 330 2282
rect 566 2278 570 2282
rect 742 2278 746 2282
rect 990 2278 994 2282
rect 1014 2278 1018 2282
rect 1046 2278 1050 2282
rect 1302 2278 1306 2282
rect 1414 2278 1418 2282
rect 1614 2278 1618 2282
rect 1870 2278 1874 2282
rect 1926 2278 1930 2282
rect 1974 2278 1978 2282
rect 2262 2278 2266 2282
rect 2510 2278 2514 2282
rect 2734 2278 2738 2282
rect 2822 2278 2826 2282
rect 2886 2278 2890 2282
rect 2974 2278 2978 2282
rect 3078 2278 3082 2282
rect 3278 2278 3282 2282
rect 3342 2278 3346 2282
rect 3366 2278 3370 2282
rect 3438 2278 3442 2282
rect 3462 2278 3466 2282
rect 3518 2278 3522 2282
rect 3694 2278 3698 2282
rect 30 2268 34 2272
rect 102 2268 106 2272
rect 134 2268 138 2272
rect 198 2268 202 2272
rect 245 2268 249 2272
rect 342 2268 346 2272
rect 422 2268 426 2272
rect 446 2268 450 2272
rect 462 2268 466 2272
rect 582 2268 586 2272
rect 758 2268 762 2272
rect 974 2268 978 2272
rect 1062 2268 1066 2272
rect 1078 2268 1082 2272
rect 1110 2268 1114 2272
rect 1118 2268 1122 2272
rect 1150 2268 1154 2272
rect 1174 2268 1178 2272
rect 1318 2268 1322 2272
rect 1406 2268 1410 2272
rect 1446 2268 1450 2272
rect 22 2258 26 2262
rect 102 2258 106 2262
rect 110 2258 114 2262
rect 206 2258 210 2262
rect 238 2258 242 2262
rect 382 2258 386 2262
rect 526 2258 530 2262
rect 702 2258 706 2262
rect 854 2258 858 2262
rect 902 2258 906 2262
rect 910 2258 914 2262
rect 950 2258 954 2262
rect 958 2258 962 2262
rect 966 2258 970 2262
rect 982 2258 986 2262
rect 998 2258 1002 2262
rect 1070 2258 1074 2262
rect 1078 2258 1082 2262
rect 1102 2258 1106 2262
rect 1134 2258 1138 2262
rect 1198 2258 1202 2262
rect 1366 2258 1370 2262
rect 1422 2258 1426 2262
rect 1446 2258 1450 2262
rect 1502 2268 1506 2272
rect 1510 2268 1514 2272
rect 1533 2268 1537 2272
rect 1630 2268 1634 2272
rect 1734 2268 1738 2272
rect 1750 2268 1754 2272
rect 1782 2268 1786 2272
rect 1790 2268 1794 2272
rect 1814 2268 1818 2272
rect 1838 2268 1842 2272
rect 1862 2268 1866 2272
rect 1902 2268 1906 2272
rect 1918 2268 1922 2272
rect 1942 2268 1946 2272
rect 1958 2268 1962 2272
rect 2030 2268 2034 2272
rect 2118 2268 2122 2272
rect 2134 2268 2138 2272
rect 2174 2268 2178 2272
rect 2278 2268 2282 2272
rect 2358 2268 2362 2272
rect 2374 2268 2378 2272
rect 2422 2268 2426 2272
rect 2454 2268 2458 2272
rect 2462 2268 2466 2272
rect 2502 2268 2506 2272
rect 2550 2268 2554 2272
rect 2582 2268 2586 2272
rect 2614 2268 2618 2272
rect 2646 2268 2650 2272
rect 2718 2268 2722 2272
rect 2830 2268 2834 2272
rect 2934 2268 2938 2272
rect 2990 2268 2994 2272
rect 3030 2268 3034 2272
rect 3038 2268 3042 2272
rect 3054 2268 3058 2272
rect 3062 2268 3066 2272
rect 3110 2268 3114 2272
rect 3150 2268 3154 2272
rect 3174 2268 3178 2272
rect 3206 2268 3210 2272
rect 3222 2268 3226 2272
rect 3270 2268 3274 2272
rect 3302 2268 3306 2272
rect 3358 2268 3362 2272
rect 3454 2268 3458 2272
rect 3486 2268 3490 2272
rect 3542 2268 3546 2272
rect 3574 2268 3578 2272
rect 1494 2258 1498 2262
rect 1574 2258 1578 2262
rect 1774 2258 1778 2262
rect 1870 2258 1874 2262
rect 1886 2258 1890 2262
rect 1950 2258 1954 2262
rect 1998 2258 2002 2262
rect 2022 2258 2026 2262
rect 2062 2258 2066 2262
rect 2094 2258 2098 2262
rect 2102 2258 2106 2262
rect 2222 2258 2226 2262
rect 2326 2258 2330 2262
rect 2366 2258 2370 2262
rect 2414 2258 2418 2262
rect 2446 2258 2450 2262
rect 2470 2258 2474 2262
rect 2486 2258 2490 2262
rect 2494 2258 2498 2262
rect 2542 2258 2546 2262
rect 2574 2258 2578 2262
rect 2606 2258 2610 2262
rect 2622 2258 2626 2262
rect 2638 2258 2642 2262
rect 2670 2258 2674 2262
rect 2774 2258 2778 2262
rect 2854 2258 2858 2262
rect 2878 2258 2882 2262
rect 2902 2258 2906 2262
rect 2966 2258 2970 2262
rect 2982 2258 2986 2262
rect 2998 2258 3002 2262
rect 3022 2258 3026 2262
rect 3038 2258 3042 2262
rect 3054 2258 3058 2262
rect 3110 2258 3114 2262
rect 3126 2258 3130 2262
rect 3150 2258 3154 2262
rect 3166 2258 3170 2262
rect 3214 2258 3218 2262
rect 3246 2258 3250 2262
rect 3302 2258 3306 2262
rect 3334 2258 3338 2262
rect 3358 2258 3362 2262
rect 3390 2258 3394 2262
rect 3398 2258 3402 2262
rect 3454 2258 3458 2262
rect 3478 2258 3482 2262
rect 3486 2258 3490 2262
rect 3518 2258 3522 2262
rect 3526 2258 3530 2262
rect 3534 2258 3538 2262
rect 3550 2258 3554 2262
rect 3614 2258 3618 2262
rect 3646 2258 3650 2262
rect 3678 2258 3682 2262
rect 3710 2258 3714 2262
rect 3734 2258 3738 2262
rect 3774 2258 3778 2262
rect 110 2248 114 2252
rect 126 2248 130 2252
rect 390 2248 394 2252
rect 470 2248 474 2252
rect 614 2250 618 2254
rect 638 2248 642 2252
rect 790 2250 794 2254
rect 1182 2248 1186 2252
rect 1350 2250 1354 2254
rect 1422 2248 1426 2252
rect 1478 2248 1482 2252
rect 1662 2250 1666 2254
rect 1702 2248 1706 2252
rect 1734 2248 1738 2252
rect 1758 2248 1762 2252
rect 1774 2248 1778 2252
rect 1790 2248 1794 2252
rect 1822 2248 1826 2252
rect 1846 2248 1850 2252
rect 2006 2248 2010 2252
rect 2310 2250 2314 2254
rect 2350 2248 2354 2252
rect 2398 2248 2402 2252
rect 2430 2248 2434 2252
rect 2486 2248 2490 2252
rect 2526 2248 2530 2252
rect 2622 2248 2626 2252
rect 2686 2250 2690 2254
rect 3006 2248 3010 2252
rect 3102 2248 3106 2252
rect 3118 2248 3122 2252
rect 3190 2248 3194 2252
rect 3254 2248 3258 2252
rect 3430 2248 3434 2252
rect 3510 2248 3514 2252
rect 3566 2248 3570 2252
rect 3590 2248 3594 2252
rect 3622 2248 3626 2252
rect 3654 2248 3658 2252
rect 3686 2248 3690 2252
rect 3742 2248 3746 2252
rect 3758 2248 3762 2252
rect 6 2238 10 2242
rect 1198 2238 1202 2242
rect 2046 2238 2050 2242
rect 2446 2238 2450 2242
rect 3134 2238 3138 2242
rect 3478 2238 3482 2242
rect 3606 2238 3610 2242
rect 3638 2238 3642 2242
rect 3670 2238 3674 2242
rect 3726 2238 3730 2242
rect 614 2227 618 2231
rect 790 2227 794 2231
rect 1350 2227 1354 2231
rect 1662 2227 1666 2231
rect 2310 2227 2314 2231
rect 2686 2227 2690 2231
rect 86 2218 90 2222
rect 390 2218 394 2222
rect 438 2218 442 2222
rect 662 2218 666 2222
rect 838 2218 842 2222
rect 886 2218 890 2222
rect 1126 2218 1130 2222
rect 1518 2218 1522 2222
rect 1966 2218 1970 2222
rect 2158 2218 2162 2222
rect 2814 2218 2818 2222
rect 2910 2218 2914 2222
rect 3126 2218 3130 2222
rect 3278 2218 3282 2222
rect 3398 2218 3402 2222
rect 3582 2218 3586 2222
rect 3614 2218 3618 2222
rect 3646 2218 3650 2222
rect 3678 2218 3682 2222
rect 3702 2218 3706 2222
rect 3734 2218 3738 2222
rect 346 2203 350 2207
rect 353 2203 357 2207
rect 1362 2203 1366 2207
rect 1369 2203 1373 2207
rect 2386 2203 2390 2207
rect 2393 2203 2397 2207
rect 3410 2203 3414 2207
rect 3417 2203 3421 2207
rect 38 2188 42 2192
rect 182 2188 186 2192
rect 478 2188 482 2192
rect 590 2188 594 2192
rect 622 2188 626 2192
rect 758 2188 762 2192
rect 862 2188 866 2192
rect 1086 2188 1090 2192
rect 1134 2188 1138 2192
rect 1214 2188 1218 2192
rect 1358 2188 1362 2192
rect 1382 2188 1386 2192
rect 1526 2188 1530 2192
rect 2014 2188 2018 2192
rect 2294 2188 2298 2192
rect 2462 2188 2466 2192
rect 2494 2188 2498 2192
rect 2558 2188 2562 2192
rect 2582 2188 2586 2192
rect 2622 2188 2626 2192
rect 2870 2188 2874 2192
rect 3014 2188 3018 2192
rect 3038 2188 3042 2192
rect 3070 2188 3074 2192
rect 3150 2188 3154 2192
rect 3510 2188 3514 2192
rect 3542 2188 3546 2192
rect 3662 2188 3666 2192
rect 3694 2188 3698 2192
rect 326 2179 330 2183
rect 558 2168 562 2172
rect 598 2168 602 2172
rect 630 2168 634 2172
rect 718 2168 722 2172
rect 782 2168 786 2172
rect 990 2179 994 2183
rect 1438 2178 1442 2182
rect 2142 2179 2146 2183
rect 3566 2168 3570 2172
rect 3598 2168 3602 2172
rect 3734 2168 3738 2172
rect 182 2158 186 2162
rect 326 2156 330 2160
rect 526 2158 530 2162
rect 574 2158 578 2162
rect 582 2158 586 2162
rect 614 2158 618 2162
rect 734 2158 738 2162
rect 798 2158 802 2162
rect 990 2156 994 2160
rect 1126 2158 1130 2162
rect 1150 2158 1154 2162
rect 1358 2158 1362 2162
rect 1494 2158 1498 2162
rect 1510 2158 1514 2162
rect 30 2148 34 2152
rect 166 2148 170 2152
rect 414 2148 418 2152
rect 494 2148 498 2152
rect 566 2148 570 2152
rect 590 2148 594 2152
rect 622 2148 626 2152
rect 678 2148 682 2152
rect 726 2148 730 2152
rect 758 2148 762 2152
rect 790 2148 794 2152
rect 822 2148 826 2152
rect 1006 2148 1010 2152
rect 1110 2148 1114 2152
rect 1126 2148 1130 2152
rect 1166 2148 1170 2152
rect 1190 2148 1194 2152
rect 1254 2148 1258 2152
rect 1454 2148 1458 2152
rect 1550 2158 1554 2162
rect 1622 2158 1626 2162
rect 1646 2158 1650 2162
rect 1662 2158 1666 2162
rect 1566 2148 1570 2152
rect 1606 2148 1610 2152
rect 1630 2148 1634 2152
rect 1702 2158 1706 2162
rect 1734 2158 1738 2162
rect 1822 2158 1826 2162
rect 1758 2148 1762 2152
rect 1790 2148 1794 2152
rect 1806 2148 1810 2152
rect 1918 2158 1922 2162
rect 1934 2158 1938 2162
rect 1950 2158 1954 2162
rect 1966 2158 1970 2162
rect 1974 2158 1978 2162
rect 2142 2156 2146 2160
rect 2214 2158 2218 2162
rect 2278 2158 2282 2162
rect 2342 2158 2346 2162
rect 2374 2158 2378 2162
rect 2390 2158 2394 2162
rect 2446 2158 2450 2162
rect 2478 2158 2482 2162
rect 2510 2158 2514 2162
rect 2518 2158 2522 2162
rect 2638 2158 2642 2162
rect 2670 2158 2674 2162
rect 2702 2158 2706 2162
rect 2718 2158 2722 2162
rect 2758 2158 2762 2162
rect 2806 2158 2810 2162
rect 1846 2148 1850 2152
rect 1918 2148 1922 2152
rect 1950 2148 1954 2152
rect 1974 2148 1978 2152
rect 1990 2148 1994 2152
rect 2158 2148 2162 2152
rect 2182 2148 2186 2152
rect 2198 2148 2202 2152
rect 2230 2148 2234 2152
rect 2246 2148 2250 2152
rect 2294 2148 2298 2152
rect 2310 2148 2314 2152
rect 2342 2148 2346 2152
rect 2358 2148 2362 2152
rect 2390 2148 2394 2152
rect 2398 2148 2402 2152
rect 2462 2148 2466 2152
rect 2494 2148 2498 2152
rect 2534 2148 2538 2152
rect 2566 2148 2570 2152
rect 2606 2148 2610 2152
rect 2662 2148 2666 2152
rect 2686 2148 2690 2152
rect 2718 2148 2722 2152
rect 2726 2148 2730 2152
rect 2750 2148 2754 2152
rect 2790 2148 2794 2152
rect 3014 2158 3018 2162
rect 3118 2158 3122 2162
rect 3198 2158 3202 2162
rect 3246 2158 3250 2162
rect 3294 2158 3298 2162
rect 3390 2158 3394 2162
rect 3526 2158 3530 2162
rect 3582 2158 3586 2162
rect 3614 2158 3618 2162
rect 3710 2158 3714 2162
rect 3718 2158 3722 2162
rect 2830 2148 2834 2152
rect 2910 2148 2914 2152
rect 3022 2148 3026 2152
rect 3110 2148 3114 2152
rect 3126 2148 3130 2152
rect 3158 2148 3162 2152
rect 3214 2148 3218 2152
rect 3254 2148 3258 2152
rect 3270 2148 3274 2152
rect 3286 2148 3290 2152
rect 3326 2148 3330 2152
rect 3342 2148 3346 2152
rect 3374 2148 3378 2152
rect 3406 2148 3410 2152
rect 3446 2148 3450 2152
rect 3470 2148 3474 2152
rect 3494 2148 3498 2152
rect 3510 2148 3514 2152
rect 3550 2148 3554 2152
rect 3574 2148 3578 2152
rect 3590 2148 3594 2152
rect 3598 2148 3602 2152
rect 3646 2148 3650 2152
rect 3678 2148 3682 2152
rect 3694 2148 3698 2152
rect 3726 2148 3730 2152
rect 3774 2148 3778 2152
rect 6 2138 10 2142
rect 134 2138 138 2142
rect 206 2138 210 2142
rect 358 2138 362 2142
rect 462 2138 466 2142
rect 502 2138 506 2142
rect 518 2138 522 2142
rect 766 2138 770 2142
rect 830 2138 834 2142
rect 958 2138 962 2142
rect 1030 2138 1034 2142
rect 1102 2138 1106 2142
rect 1166 2138 1170 2142
rect 1198 2138 1202 2142
rect 1310 2138 1314 2142
rect 1446 2138 1450 2142
rect 1462 2138 1466 2142
rect 1486 2138 1490 2142
rect 1494 2138 1498 2142
rect 1518 2138 1522 2142
rect 1630 2138 1634 2142
rect 1646 2138 1650 2142
rect 1670 2138 1674 2142
rect 1694 2138 1698 2142
rect 1726 2138 1730 2142
rect 1766 2138 1770 2142
rect 1774 2138 1778 2142
rect 1798 2138 1802 2142
rect 1838 2138 1842 2142
rect 1878 2138 1882 2142
rect 1910 2138 1914 2142
rect 1942 2138 1946 2142
rect 1998 2138 2002 2142
rect 2110 2138 2114 2142
rect 2206 2138 2210 2142
rect 2222 2138 2226 2142
rect 2238 2138 2242 2142
rect 2254 2138 2258 2142
rect 2302 2138 2306 2142
rect 2318 2138 2322 2142
rect 2366 2138 2370 2142
rect 2414 2138 2418 2142
rect 2422 2138 2426 2142
rect 2438 2138 2442 2142
rect 2454 2138 2458 2142
rect 2486 2138 2490 2142
rect 2550 2138 2554 2142
rect 2662 2138 2666 2142
rect 2694 2138 2698 2142
rect 2726 2138 2730 2142
rect 2734 2138 2738 2142
rect 2774 2138 2778 2142
rect 2782 2138 2786 2142
rect 2822 2138 2826 2142
rect 2838 2138 2842 2142
rect 2966 2138 2970 2142
rect 3054 2138 3058 2142
rect 3086 2138 3090 2142
rect 3102 2138 3106 2142
rect 3134 2138 3138 2142
rect 3150 2138 3154 2142
rect 3182 2138 3186 2142
rect 3222 2138 3226 2142
rect 3230 2138 3234 2142
rect 3246 2138 3250 2142
rect 3278 2138 3282 2142
rect 3294 2138 3298 2142
rect 3310 2138 3314 2142
rect 3334 2138 3338 2142
rect 3566 2138 3570 2142
rect 3686 2138 3690 2142
rect 118 2128 122 2132
rect 374 2128 378 2132
rect 454 2128 458 2132
rect 942 2128 946 2132
rect 1142 2128 1146 2132
rect 1294 2128 1298 2132
rect 1406 2128 1410 2132
rect 1582 2128 1586 2132
rect 1862 2128 1866 2132
rect 2094 2128 2098 2132
rect 2270 2128 2274 2132
rect 2334 2128 2338 2132
rect 2342 2128 2346 2132
rect 2550 2128 2554 2132
rect 2766 2128 2770 2132
rect 2950 2128 2954 2132
rect 3062 2128 3066 2132
rect 3094 2128 3098 2132
rect 3150 2128 3154 2132
rect 3182 2128 3186 2132
rect 3318 2128 3322 2132
rect 3430 2128 3434 2132
rect 3470 2128 3474 2132
rect 3478 2128 3482 2132
rect 3534 2128 3538 2132
rect 262 2118 266 2122
rect 478 2118 482 2122
rect 510 2118 514 2122
rect 654 2118 658 2122
rect 694 2118 698 2122
rect 806 2118 810 2122
rect 1478 2118 1482 2122
rect 2262 2118 2266 2122
rect 2518 2118 2522 2122
rect 2582 2118 2586 2122
rect 2638 2118 2642 2122
rect 2670 2118 2674 2122
rect 3246 2118 3250 2122
rect 3438 2118 3442 2122
rect 3630 2118 3634 2122
rect 3742 2118 3746 2122
rect 3758 2118 3762 2122
rect 850 2103 854 2107
rect 857 2103 861 2107
rect 1882 2103 1886 2107
rect 1889 2103 1893 2107
rect 2906 2103 2910 2107
rect 2913 2103 2917 2107
rect 638 2088 642 2092
rect 646 2088 650 2092
rect 1126 2088 1130 2092
rect 1158 2088 1162 2092
rect 1198 2088 1202 2092
rect 1278 2088 1282 2092
rect 1310 2088 1314 2092
rect 1518 2088 1522 2092
rect 1718 2088 1722 2092
rect 1846 2088 1850 2092
rect 1870 2088 1874 2092
rect 1974 2088 1978 2092
rect 2230 2088 2234 2092
rect 2278 2088 2282 2092
rect 2294 2088 2298 2092
rect 2342 2088 2346 2092
rect 2470 2088 2474 2092
rect 2502 2088 2506 2092
rect 2558 2088 2562 2092
rect 2646 2088 2650 2092
rect 2734 2088 2738 2092
rect 2990 2088 2994 2092
rect 3046 2088 3050 2092
rect 3142 2088 3146 2092
rect 3174 2088 3178 2092
rect 3206 2088 3210 2092
rect 3278 2088 3282 2092
rect 3574 2088 3578 2092
rect 3598 2088 3602 2092
rect 3654 2088 3658 2092
rect 3678 2088 3682 2092
rect 206 2078 210 2082
rect 398 2078 402 2082
rect 598 2078 602 2082
rect 758 2078 762 2082
rect 1046 2078 1050 2082
rect 1222 2078 1226 2082
rect 1238 2078 1242 2082
rect 1406 2078 1410 2082
rect 1470 2078 1474 2082
rect 6 2068 10 2072
rect 30 2068 34 2072
rect 54 2068 58 2072
rect 86 2068 90 2072
rect 222 2068 226 2072
rect 414 2068 418 2072
rect 486 2068 490 2072
rect 502 2068 506 2072
rect 518 2068 522 2072
rect 566 2068 570 2072
rect 582 2068 586 2072
rect 670 2068 674 2072
rect 742 2068 746 2072
rect 870 2068 874 2072
rect 1030 2068 1034 2072
rect 1214 2068 1218 2072
rect 1246 2068 1250 2072
rect 1366 2068 1370 2072
rect 1422 2068 1426 2072
rect 1470 2068 1474 2072
rect 1486 2068 1490 2072
rect 1510 2068 1514 2072
rect 1534 2078 1538 2082
rect 1638 2078 1642 2082
rect 1838 2078 1842 2082
rect 1862 2078 1866 2082
rect 1902 2078 1906 2082
rect 1942 2078 1946 2082
rect 2054 2078 2058 2082
rect 2286 2078 2290 2082
rect 2310 2078 2314 2082
rect 2350 2078 2354 2082
rect 2534 2078 2538 2082
rect 2566 2078 2570 2082
rect 2686 2078 2690 2082
rect 2822 2078 2826 2082
rect 2966 2078 2970 2082
rect 3038 2078 3042 2082
rect 3054 2078 3058 2082
rect 3094 2078 3098 2082
rect 3150 2078 3154 2082
rect 3182 2078 3186 2082
rect 3214 2078 3218 2082
rect 3222 2078 3226 2082
rect 3246 2078 3250 2082
rect 3294 2078 3298 2082
rect 3342 2078 3346 2082
rect 3366 2078 3370 2082
rect 3470 2078 3474 2082
rect 3646 2078 3650 2082
rect 3766 2078 3770 2082
rect 1622 2068 1626 2072
rect 1726 2068 1730 2072
rect 1766 2068 1770 2072
rect 1782 2068 1786 2072
rect 1830 2068 1834 2072
rect 1878 2068 1882 2072
rect 2070 2068 2074 2072
rect 2150 2068 2154 2072
rect 22 2058 26 2062
rect 54 2058 58 2062
rect 62 2058 66 2062
rect 94 2058 98 2062
rect 166 2058 170 2062
rect 222 2058 226 2062
rect 270 2058 274 2062
rect 317 2058 321 2062
rect 358 2058 362 2062
rect 462 2058 466 2062
rect 510 2058 514 2062
rect 542 2058 546 2062
rect 574 2058 578 2062
rect 622 2058 626 2062
rect 670 2058 674 2062
rect 702 2058 706 2062
rect 798 2058 802 2062
rect 878 2058 882 2062
rect 894 2058 898 2062
rect 918 2058 922 2062
rect 950 2058 954 2062
rect 982 2058 986 2062
rect 1150 2058 1154 2062
rect 1182 2058 1186 2062
rect 1238 2058 1242 2062
rect 1262 2058 1266 2062
rect 1294 2058 1298 2062
rect 1390 2058 1394 2062
rect 1446 2058 1450 2062
rect 1462 2058 1466 2062
rect 1494 2058 1498 2062
rect 1502 2058 1506 2062
rect 1550 2058 1554 2062
rect 1582 2058 1586 2062
rect 1742 2058 1746 2062
rect 1822 2058 1826 2062
rect 1854 2058 1858 2062
rect 1886 2058 1890 2062
rect 1926 2058 1930 2062
rect 1934 2058 1938 2062
rect 1958 2058 1962 2062
rect 2014 2058 2018 2062
rect 2070 2058 2074 2062
rect 2190 2068 2194 2072
rect 2222 2068 2226 2072
rect 2270 2068 2274 2072
rect 2302 2068 2306 2072
rect 2326 2068 2330 2072
rect 2390 2068 2394 2072
rect 2414 2068 2418 2072
rect 2542 2068 2546 2072
rect 2550 2068 2554 2072
rect 2566 2068 2570 2072
rect 2590 2068 2594 2072
rect 2606 2068 2610 2072
rect 2654 2068 2658 2072
rect 2718 2068 2722 2072
rect 2726 2068 2730 2072
rect 2806 2068 2810 2072
rect 2950 2068 2954 2072
rect 2982 2068 2986 2072
rect 3030 2068 3034 2072
rect 3118 2068 3122 2072
rect 3134 2068 3138 2072
rect 3166 2068 3170 2072
rect 3198 2068 3202 2072
rect 3294 2068 3298 2072
rect 3302 2068 3306 2072
rect 3318 2068 3322 2072
rect 3390 2068 3394 2072
rect 3438 2068 3442 2072
rect 3606 2068 3610 2072
rect 3710 2068 3714 2072
rect 2166 2058 2170 2062
rect 2206 2058 2210 2062
rect 2262 2058 2266 2062
rect 2310 2058 2314 2062
rect 2326 2058 2330 2062
rect 2366 2058 2370 2062
rect 2398 2058 2402 2062
rect 2422 2058 2426 2062
rect 2454 2058 2458 2062
rect 2486 2058 2490 2062
rect 2518 2058 2522 2062
rect 2582 2058 2586 2062
rect 2614 2058 2618 2062
rect 2662 2058 2666 2062
rect 2670 2058 2674 2062
rect 2710 2058 2714 2062
rect 2806 2058 2810 2062
rect 2862 2058 2866 2062
rect 2950 2058 2954 2062
rect 2974 2058 2978 2062
rect 3022 2058 3026 2062
rect 3054 2058 3058 2062
rect 3086 2058 3090 2062
rect 3118 2058 3122 2062
rect 3126 2058 3130 2062
rect 3158 2058 3162 2062
rect 3190 2058 3194 2062
rect 3222 2058 3226 2062
rect 3238 2058 3242 2062
rect 3262 2058 3266 2062
rect 3310 2058 3314 2062
rect 3358 2058 3362 2062
rect 3382 2058 3386 2062
rect 3398 2058 3402 2062
rect 3446 2058 3450 2062
rect 3470 2058 3474 2062
rect 3486 2058 3490 2062
rect 3502 2058 3506 2062
rect 3542 2058 3546 2062
rect 3574 2058 3578 2062
rect 3622 2058 3626 2062
rect 3662 2058 3666 2062
rect 3678 2058 3682 2062
rect 3718 2058 3722 2062
rect 3742 2058 3746 2062
rect 62 2048 66 2052
rect 78 2048 82 2052
rect 254 2050 258 2054
rect 446 2050 450 2054
rect 526 2048 530 2052
rect 534 2048 538 2052
rect 590 2048 594 2052
rect 646 2048 650 2052
rect 710 2050 714 2054
rect 926 2048 930 2052
rect 958 2048 962 2052
rect 998 2050 1002 2054
rect 1142 2048 1146 2052
rect 1174 2048 1178 2052
rect 1462 2048 1466 2052
rect 1590 2050 1594 2054
rect 1758 2048 1762 2052
rect 1806 2048 1810 2052
rect 1910 2048 1914 2052
rect 2102 2050 2106 2054
rect 2182 2048 2186 2052
rect 2214 2048 2218 2052
rect 2446 2048 2450 2052
rect 2502 2048 2506 2052
rect 2598 2048 2602 2052
rect 2630 2048 2634 2052
rect 2694 2048 2698 2052
rect 2758 2048 2762 2052
rect 3006 2048 3010 2052
rect 3270 2048 3274 2052
rect 3334 2048 3338 2052
rect 3414 2048 3418 2052
rect 3462 2048 3466 2052
rect 3518 2048 3522 2052
rect 3550 2048 3554 2052
rect 3582 2048 3586 2052
rect 3590 2048 3594 2052
rect 3638 2048 3642 2052
rect 3670 2048 3674 2052
rect 3726 2048 3730 2052
rect 3734 2048 3738 2052
rect 94 2038 98 2042
rect 550 2038 554 2042
rect 862 2038 866 2042
rect 910 2038 914 2042
rect 942 2038 946 2042
rect 1158 2038 1162 2042
rect 1190 2038 1194 2042
rect 1206 2038 1210 2042
rect 1742 2038 1746 2042
rect 1782 2038 1786 2042
rect 2374 2038 2378 2042
rect 2678 2038 2682 2042
rect 3358 2038 3362 2042
rect 3382 2038 3386 2042
rect 3502 2038 3506 2042
rect 3534 2038 3538 2042
rect 3566 2038 3570 2042
rect 3622 2038 3626 2042
rect 3686 2038 3690 2042
rect 3718 2038 3722 2042
rect 3750 2038 3754 2042
rect 446 2027 450 2031
rect 998 2027 1002 2031
rect 1590 2027 1594 2031
rect 2102 2027 2106 2031
rect 2430 2028 2434 2032
rect 2902 2028 2906 2032
rect 3742 2028 3746 2032
rect 126 2018 130 2022
rect 254 2018 258 2022
rect 542 2018 546 2022
rect 710 2018 714 2022
rect 950 2018 954 2022
rect 1198 2018 1202 2022
rect 1230 2018 1234 2022
rect 1254 2018 1258 2022
rect 1406 2018 1410 2022
rect 1430 2018 1434 2022
rect 1774 2018 1778 2022
rect 2142 2018 2146 2022
rect 2230 2018 2234 2022
rect 2294 2018 2298 2022
rect 2758 2018 2762 2022
rect 3094 2018 3098 2022
rect 3262 2018 3266 2022
rect 3326 2018 3330 2022
rect 3398 2018 3402 2022
rect 3542 2018 3546 2022
rect 3630 2018 3634 2022
rect 3774 2018 3778 2022
rect 346 2003 350 2007
rect 353 2003 357 2007
rect 1362 2003 1366 2007
rect 1369 2003 1373 2007
rect 2386 2003 2390 2007
rect 2393 2003 2397 2007
rect 3410 2003 3414 2007
rect 3417 2003 3421 2007
rect 6 1988 10 1992
rect 238 1988 242 1992
rect 270 1988 274 1992
rect 526 1988 530 1992
rect 590 1988 594 1992
rect 654 1988 658 1992
rect 710 1988 714 1992
rect 878 1988 882 1992
rect 950 1988 954 1992
rect 1014 1988 1018 1992
rect 1030 1988 1034 1992
rect 1070 1988 1074 1992
rect 1126 1988 1130 1992
rect 1166 1988 1170 1992
rect 1182 1988 1186 1992
rect 1214 1988 1218 1992
rect 1358 1988 1362 1992
rect 1470 1988 1474 1992
rect 1542 1988 1546 1992
rect 1566 1988 1570 1992
rect 1726 1988 1730 1992
rect 1790 1988 1794 1992
rect 1862 1988 1866 1992
rect 1974 1988 1978 1992
rect 2030 1988 2034 1992
rect 2174 1988 2178 1992
rect 2470 1988 2474 1992
rect 2830 1988 2834 1992
rect 2854 1988 2858 1992
rect 2942 1988 2946 1992
rect 3014 1988 3018 1992
rect 3718 1988 3722 1992
rect 30 1968 34 1972
rect 382 1968 386 1972
rect 1630 1978 1634 1982
rect 2326 1978 2330 1982
rect 630 1968 634 1972
rect 662 1968 666 1972
rect 1062 1968 1066 1972
rect 1078 1968 1082 1972
rect 1102 1968 1106 1972
rect 1134 1968 1138 1972
rect 1158 1968 1162 1972
rect 1166 1968 1170 1972
rect 1478 1968 1482 1972
rect 1758 1968 1762 1972
rect 3710 1968 3714 1972
rect 3726 1968 3730 1972
rect 62 1958 66 1962
rect 238 1958 242 1962
rect 286 1958 290 1962
rect 526 1958 530 1962
rect 550 1958 554 1962
rect 614 1958 618 1962
rect 646 1958 650 1962
rect 678 1958 682 1962
rect 878 1958 882 1962
rect 918 1958 922 1962
rect 998 1958 1002 1962
rect 1118 1958 1122 1962
rect 1174 1958 1178 1962
rect 1214 1958 1218 1962
rect 22 1948 26 1952
rect 46 1948 50 1952
rect 62 1948 66 1952
rect 222 1948 226 1952
rect 262 1948 266 1952
rect 310 1948 314 1952
rect 334 1948 338 1952
rect 478 1948 482 1952
rect 550 1948 554 1952
rect 566 1948 570 1952
rect 590 1948 594 1952
rect 622 1948 626 1952
rect 662 1948 666 1952
rect 678 1948 682 1952
rect 694 1948 698 1952
rect 726 1948 730 1952
rect 774 1948 778 1952
rect 926 1948 930 1952
rect 934 1948 938 1952
rect 990 1948 994 1952
rect 1014 1948 1018 1952
rect 1046 1948 1050 1952
rect 1054 1948 1058 1952
rect 1070 1948 1074 1952
rect 1126 1948 1130 1952
rect 1158 1948 1162 1952
rect 1166 1948 1170 1952
rect 1318 1948 1322 1952
rect 1430 1958 1434 1962
rect 1462 1958 1466 1962
rect 1582 1958 1586 1962
rect 1446 1948 1450 1952
rect 1470 1948 1474 1952
rect 1494 1948 1498 1952
rect 1518 1948 1522 1952
rect 1566 1948 1570 1952
rect 1590 1948 1594 1952
rect 1606 1948 1610 1952
rect 1630 1948 1634 1952
rect 1654 1958 1658 1962
rect 1710 1958 1714 1962
rect 1742 1958 1746 1962
rect 1774 1958 1778 1962
rect 1806 1958 1810 1962
rect 2174 1958 2178 1962
rect 2198 1958 2202 1962
rect 2262 1958 2266 1962
rect 2342 1958 2346 1962
rect 2430 1958 2434 1962
rect 2478 1958 2482 1962
rect 2510 1958 2514 1962
rect 2542 1958 2546 1962
rect 2598 1958 2602 1962
rect 2662 1958 2666 1962
rect 2694 1958 2698 1962
rect 2734 1958 2738 1962
rect 2750 1958 2754 1962
rect 2790 1958 2794 1962
rect 2870 1958 2874 1962
rect 2926 1958 2930 1962
rect 2958 1958 2962 1962
rect 3022 1958 3026 1962
rect 3094 1958 3098 1962
rect 3182 1958 3186 1962
rect 3382 1958 3386 1962
rect 3502 1958 3506 1962
rect 3582 1958 3586 1962
rect 3638 1958 3642 1962
rect 3726 1958 3730 1962
rect 3734 1958 3738 1962
rect 1670 1948 1674 1952
rect 1694 1948 1698 1952
rect 1726 1948 1730 1952
rect 1758 1948 1762 1952
rect 1790 1948 1794 1952
rect 1814 1948 1818 1952
rect 1830 1948 1834 1952
rect 1846 1948 1850 1952
rect 1870 1948 1874 1952
rect 1958 1948 1962 1952
rect 1990 1948 1994 1952
rect 2022 1948 2026 1952
rect 2070 1948 2074 1952
rect 2158 1948 2162 1952
rect 2198 1948 2202 1952
rect 2214 1948 2218 1952
rect 2254 1948 2258 1952
rect 2262 1948 2266 1952
rect 2278 1948 2282 1952
rect 2294 1948 2298 1952
rect 2326 1948 2330 1952
rect 2350 1948 2354 1952
rect 2366 1948 2370 1952
rect 2382 1948 2386 1952
rect 2398 1948 2402 1952
rect 2438 1948 2442 1952
rect 2446 1948 2450 1952
rect 2526 1948 2530 1952
rect 2558 1948 2562 1952
rect 2582 1948 2586 1952
rect 2710 1948 2714 1952
rect 2734 1948 2738 1952
rect 2758 1948 2762 1952
rect 2774 1948 2778 1952
rect 2814 1948 2818 1952
rect 2854 1948 2858 1952
rect 2878 1948 2882 1952
rect 2894 1948 2898 1952
rect 2942 1948 2946 1952
rect 2982 1948 2986 1952
rect 3030 1948 3034 1952
rect 3062 1948 3066 1952
rect 3078 1948 3082 1952
rect 3110 1948 3114 1952
rect 3158 1948 3162 1952
rect 3214 1948 3218 1952
rect 3238 1948 3242 1952
rect 3262 1948 3266 1952
rect 3278 1948 3282 1952
rect 3302 1948 3306 1952
rect 3310 1948 3314 1952
rect 3342 1948 3346 1952
rect 3374 1948 3378 1952
rect 3446 1948 3450 1952
rect 3478 1948 3482 1952
rect 3486 1948 3490 1952
rect 3526 1948 3530 1952
rect 3550 1948 3554 1952
rect 3566 1948 3570 1952
rect 3606 1948 3610 1952
rect 3630 1948 3634 1952
rect 3654 1948 3658 1952
rect 3694 1948 3698 1952
rect 3718 1948 3722 1952
rect 3742 1948 3746 1952
rect 54 1938 58 1942
rect 190 1938 194 1942
rect 262 1938 266 1942
rect 294 1938 298 1942
rect 358 1938 362 1942
rect 478 1938 482 1942
rect 574 1938 578 1942
rect 582 1938 586 1942
rect 702 1938 706 1942
rect 830 1938 834 1942
rect 1022 1938 1026 1942
rect 1094 1938 1098 1942
rect 1190 1938 1194 1942
rect 1262 1938 1266 1942
rect 1398 1938 1402 1942
rect 1406 1938 1410 1942
rect 1454 1938 1458 1942
rect 1558 1938 1562 1942
rect 1590 1938 1594 1942
rect 1622 1938 1626 1942
rect 1678 1938 1682 1942
rect 1686 1938 1690 1942
rect 1718 1938 1722 1942
rect 1750 1938 1754 1942
rect 1782 1938 1786 1942
rect 1822 1938 1826 1942
rect 1934 1938 1938 1942
rect 1990 1938 1994 1942
rect 2126 1938 2130 1942
rect 2246 1938 2250 1942
rect 2286 1938 2290 1942
rect 2318 1938 2322 1942
rect 2350 1938 2354 1942
rect 2406 1938 2410 1942
rect 2454 1938 2458 1942
rect 2462 1938 2466 1942
rect 2486 1938 2490 1942
rect 2502 1938 2506 1942
rect 2534 1938 2538 1942
rect 2566 1938 2570 1942
rect 2574 1938 2578 1942
rect 2598 1938 2602 1942
rect 2646 1938 2650 1942
rect 2686 1938 2690 1942
rect 2718 1938 2722 1942
rect 2726 1938 2730 1942
rect 2766 1938 2770 1942
rect 2806 1938 2810 1942
rect 2846 1938 2850 1942
rect 2886 1938 2890 1942
rect 2950 1938 2954 1942
rect 2974 1938 2978 1942
rect 2998 1938 3002 1942
rect 3006 1938 3010 1942
rect 3022 1938 3026 1942
rect 3038 1938 3042 1942
rect 3054 1938 3058 1942
rect 3070 1938 3074 1942
rect 3102 1938 3106 1942
rect 3150 1938 3154 1942
rect 3166 1938 3170 1942
rect 3206 1938 3210 1942
rect 3310 1938 3314 1942
rect 3398 1938 3402 1942
rect 3414 1938 3418 1942
rect 3438 1938 3442 1942
rect 3454 1938 3458 1942
rect 3470 1938 3474 1942
rect 3526 1938 3530 1942
rect 3558 1938 3562 1942
rect 174 1928 178 1932
rect 462 1928 466 1932
rect 718 1928 722 1932
rect 814 1928 818 1932
rect 958 1928 962 1932
rect 1278 1928 1282 1932
rect 1510 1928 1514 1932
rect 1534 1928 1538 1932
rect 1550 1928 1554 1932
rect 1614 1928 1618 1932
rect 1838 1928 1842 1932
rect 1910 1928 1914 1932
rect 1926 1928 1930 1932
rect 2110 1928 2114 1932
rect 2230 1928 2234 1932
rect 2310 1928 2314 1932
rect 2382 1928 2386 1932
rect 2422 1928 2426 1932
rect 2622 1928 2626 1932
rect 2782 1928 2786 1932
rect 2798 1928 2802 1932
rect 2902 1928 2906 1932
rect 2958 1928 2962 1932
rect 2990 1928 2994 1932
rect 3134 1928 3138 1932
rect 3190 1928 3194 1932
rect 3222 1928 3226 1932
rect 3254 1928 3258 1932
rect 3278 1928 3282 1932
rect 3286 1928 3290 1932
rect 3302 1928 3306 1932
rect 3334 1928 3338 1932
rect 3422 1928 3426 1932
rect 3454 1928 3458 1932
rect 3510 1928 3514 1932
rect 3630 1938 3634 1942
rect 3662 1938 3666 1942
rect 3670 1938 3674 1942
rect 3534 1928 3538 1932
rect 3550 1928 3554 1932
rect 3590 1928 3594 1932
rect 3606 1928 3610 1932
rect 3614 1928 3618 1932
rect 94 1918 98 1922
rect 302 1918 306 1922
rect 366 1918 370 1922
rect 710 1918 714 1922
rect 974 1918 978 1922
rect 1038 1918 1042 1922
rect 1070 1918 1074 1922
rect 1142 1918 1146 1922
rect 1414 1918 1418 1922
rect 1502 1918 1506 1922
rect 1526 1918 1530 1922
rect 1710 1918 1714 1922
rect 1862 1918 1866 1922
rect 1950 1918 1954 1922
rect 1974 1918 1978 1922
rect 2414 1918 2418 1922
rect 2470 1918 2474 1922
rect 2542 1918 2546 1922
rect 2638 1918 2642 1922
rect 3046 1918 3050 1922
rect 3094 1918 3098 1922
rect 3126 1918 3130 1922
rect 3182 1918 3186 1922
rect 3198 1918 3202 1922
rect 3246 1918 3250 1922
rect 3366 1918 3370 1922
rect 3502 1918 3506 1922
rect 3582 1918 3586 1922
rect 3638 1918 3642 1922
rect 3742 1918 3746 1922
rect 850 1903 854 1907
rect 857 1903 861 1907
rect 1882 1903 1886 1907
rect 1889 1903 1893 1907
rect 2906 1903 2910 1907
rect 2913 1903 2917 1907
rect 30 1888 34 1892
rect 518 1888 522 1892
rect 646 1888 650 1892
rect 662 1888 666 1892
rect 702 1888 706 1892
rect 734 1888 738 1892
rect 806 1888 810 1892
rect 846 1888 850 1892
rect 1230 1888 1234 1892
rect 1318 1888 1322 1892
rect 1390 1888 1394 1892
rect 1534 1888 1538 1892
rect 1558 1888 1562 1892
rect 1590 1888 1594 1892
rect 1614 1888 1618 1892
rect 1646 1888 1650 1892
rect 1694 1888 1698 1892
rect 2294 1888 2298 1892
rect 2350 1888 2354 1892
rect 2366 1888 2370 1892
rect 2446 1888 2450 1892
rect 2478 1888 2482 1892
rect 2742 1888 2746 1892
rect 2942 1888 2946 1892
rect 2982 1888 2986 1892
rect 3014 1888 3018 1892
rect 3046 1888 3050 1892
rect 3062 1888 3066 1892
rect 3102 1888 3106 1892
rect 3206 1888 3210 1892
rect 3446 1888 3450 1892
rect 134 1878 138 1882
rect 318 1878 322 1882
rect 918 1878 922 1882
rect 926 1878 930 1882
rect 1054 1878 1058 1882
rect 1078 1878 1082 1882
rect 1198 1878 1202 1882
rect 1206 1878 1210 1882
rect 1214 1878 1218 1882
rect 1326 1878 1330 1882
rect 1574 1878 1578 1882
rect 1790 1878 1794 1882
rect 2038 1878 2042 1882
rect 2086 1878 2090 1882
rect 2190 1878 2194 1882
rect 2270 1878 2274 1882
rect 2430 1878 2434 1882
rect 150 1868 154 1872
rect 222 1868 226 1872
rect 302 1868 306 1872
rect 406 1868 410 1872
rect 462 1868 466 1872
rect 478 1868 482 1872
rect 494 1868 498 1872
rect 534 1868 538 1872
rect 550 1868 554 1872
rect 590 1868 594 1872
rect 606 1868 610 1872
rect 622 1868 626 1872
rect 654 1868 658 1872
rect 678 1868 682 1872
rect 710 1868 714 1872
rect 742 1868 746 1872
rect 790 1868 794 1872
rect 814 1868 818 1872
rect 822 1868 826 1872
rect 838 1868 842 1872
rect 862 1868 866 1872
rect 934 1868 938 1872
rect 966 1868 970 1872
rect 1030 1868 1034 1872
rect 1046 1868 1050 1872
rect 1102 1868 1106 1872
rect 1126 1868 1130 1872
rect 1158 1868 1162 1872
rect 1238 1868 1242 1872
rect 1270 1868 1274 1872
rect 1302 1868 1306 1872
rect 1334 1868 1338 1872
rect 1486 1868 1490 1872
rect 1510 1868 1514 1872
rect 1518 1868 1522 1872
rect 1542 1868 1546 1872
rect 1582 1868 1586 1872
rect 1614 1868 1618 1872
rect 1630 1868 1634 1872
rect 1670 1868 1674 1872
rect 1678 1868 1682 1872
rect 1806 1868 1810 1872
rect 1894 1868 1898 1872
rect 1926 1868 1930 1872
rect 1950 1868 1954 1872
rect 1982 1868 1986 1872
rect 2014 1868 2018 1872
rect 2030 1868 2034 1872
rect 2174 1868 2178 1872
rect 2286 1868 2290 1872
rect 2302 1868 2306 1872
rect 2318 1868 2322 1872
rect 2334 1868 2338 1872
rect 2366 1868 2370 1872
rect 2406 1868 2410 1872
rect 2662 1878 2666 1882
rect 2838 1878 2842 1882
rect 2846 1878 2850 1882
rect 2878 1878 2882 1882
rect 2918 1878 2922 1882
rect 3038 1878 3042 1882
rect 3086 1878 3090 1882
rect 3246 1878 3250 1882
rect 3254 1878 3258 1882
rect 3286 1878 3290 1882
rect 3318 1878 3322 1882
rect 3382 1878 3386 1882
rect 3454 1878 3458 1882
rect 3478 1878 3482 1882
rect 3534 1878 3538 1882
rect 3590 1878 3594 1882
rect 3606 1878 3610 1882
rect 2454 1868 2458 1872
rect 2462 1868 2466 1872
rect 2510 1868 2514 1872
rect 2518 1868 2522 1872
rect 2534 1868 2538 1872
rect 2550 1868 2554 1872
rect 2646 1868 2650 1872
rect 2758 1868 2762 1872
rect 2782 1868 2786 1872
rect 2822 1868 2826 1872
rect 2846 1868 2850 1872
rect 2934 1868 2938 1872
rect 2950 1868 2954 1872
rect 2974 1868 2978 1872
rect 2998 1868 3002 1872
rect 3078 1868 3082 1872
rect 3158 1868 3162 1872
rect 3198 1868 3202 1872
rect 3214 1868 3218 1872
rect 3270 1868 3274 1872
rect 3302 1868 3306 1872
rect 3334 1868 3338 1872
rect 3422 1868 3426 1872
rect 3470 1868 3474 1872
rect 3494 1868 3498 1872
rect 3614 1868 3618 1872
rect 198 1858 202 1862
rect 182 1850 186 1854
rect 358 1858 362 1862
rect 454 1858 458 1862
rect 470 1858 474 1862
rect 494 1858 498 1862
rect 542 1858 546 1862
rect 566 1858 570 1862
rect 598 1858 602 1862
rect 630 1858 634 1862
rect 686 1858 690 1862
rect 718 1858 722 1862
rect 782 1858 786 1862
rect 902 1858 906 1862
rect 942 1858 946 1862
rect 990 1858 994 1862
rect 1062 1858 1066 1862
rect 1102 1858 1106 1862
rect 1142 1858 1146 1862
rect 1294 1858 1298 1862
rect 1430 1858 1434 1862
rect 1510 1858 1514 1862
rect 1606 1858 1610 1862
rect 1638 1858 1642 1862
rect 1662 1858 1666 1862
rect 1854 1858 1858 1862
rect 1902 1858 1906 1862
rect 2006 1858 2010 1862
rect 2022 1858 2026 1862
rect 2070 1858 2074 1862
rect 2078 1858 2082 1862
rect 2102 1858 2106 1862
rect 2230 1858 2234 1862
rect 2310 1858 2314 1862
rect 2358 1858 2362 1862
rect 2390 1858 2394 1862
rect 2414 1858 2418 1862
rect 2470 1858 2474 1862
rect 2502 1858 2506 1862
rect 2526 1858 2530 1862
rect 2542 1858 2546 1862
rect 2606 1858 2610 1862
rect 2790 1858 2794 1862
rect 2814 1858 2818 1862
rect 2830 1858 2834 1862
rect 2870 1858 2874 1862
rect 2894 1858 2898 1862
rect 2934 1858 2938 1862
rect 3030 1858 3034 1862
rect 3054 1858 3058 1862
rect 3118 1858 3122 1862
rect 3142 1858 3146 1862
rect 3166 1858 3170 1862
rect 3182 1858 3186 1862
rect 3222 1858 3226 1862
rect 3230 1858 3234 1862
rect 3246 1858 3250 1862
rect 3278 1858 3282 1862
rect 3310 1858 3314 1862
rect 3342 1858 3346 1862
rect 3374 1858 3378 1862
rect 3398 1858 3402 1862
rect 3470 1858 3474 1862
rect 3494 1858 3498 1862
rect 3510 1858 3514 1862
rect 3550 1858 3554 1862
rect 3574 1858 3578 1862
rect 3606 1858 3610 1862
rect 3622 1858 3626 1862
rect 3638 1858 3642 1862
rect 3654 1858 3658 1862
rect 3694 1858 3698 1862
rect 3726 1858 3730 1862
rect 3758 1858 3762 1862
rect 246 1848 250 1852
rect 270 1850 274 1854
rect 486 1848 490 1852
rect 526 1848 530 1852
rect 558 1848 562 1852
rect 614 1848 618 1852
rect 646 1848 650 1852
rect 670 1848 674 1852
rect 702 1848 706 1852
rect 734 1848 738 1852
rect 758 1848 762 1852
rect 798 1848 802 1852
rect 822 1848 826 1852
rect 846 1848 850 1852
rect 910 1848 914 1852
rect 950 1848 954 1852
rect 966 1848 970 1852
rect 998 1848 1002 1852
rect 1118 1848 1122 1852
rect 1174 1848 1178 1852
rect 1222 1848 1226 1852
rect 1246 1848 1250 1852
rect 1262 1848 1266 1852
rect 1278 1848 1282 1852
rect 1422 1848 1426 1852
rect 1478 1848 1482 1852
rect 1534 1848 1538 1852
rect 1598 1848 1602 1852
rect 1646 1848 1650 1852
rect 1694 1848 1698 1852
rect 1838 1850 1842 1854
rect 1918 1848 1922 1852
rect 1958 1848 1962 1852
rect 1990 1848 1994 1852
rect 2054 1848 2058 1852
rect 2142 1850 2146 1854
rect 2326 1848 2330 1852
rect 2350 1848 2354 1852
rect 2486 1848 2490 1852
rect 2542 1848 2546 1852
rect 2574 1848 2578 1852
rect 2598 1848 2602 1852
rect 2774 1848 2778 1852
rect 2790 1848 2794 1852
rect 2806 1848 2810 1852
rect 2950 1848 2954 1852
rect 2982 1848 2986 1852
rect 3150 1848 3154 1852
rect 3166 1848 3170 1852
rect 3182 1848 3186 1852
rect 3254 1848 3258 1852
rect 3446 1848 3450 1852
rect 3526 1848 3530 1852
rect 3582 1848 3586 1852
rect 3638 1848 3642 1852
rect 3670 1848 3674 1852
rect 3702 1848 3706 1852
rect 3734 1848 3738 1852
rect 3766 1848 3770 1852
rect 566 1838 570 1842
rect 574 1838 578 1842
rect 654 1838 658 1842
rect 894 1838 898 1842
rect 982 1838 986 1842
rect 1438 1838 1442 1842
rect 1558 1838 1562 1842
rect 3134 1838 3138 1842
rect 3494 1838 3498 1842
rect 3566 1838 3570 1842
rect 3662 1838 3666 1842
rect 3686 1838 3690 1842
rect 3718 1838 3722 1842
rect 3750 1838 3754 1842
rect 270 1827 274 1831
rect 2142 1827 2146 1831
rect 3286 1828 3290 1832
rect 3550 1828 3554 1832
rect 182 1818 186 1822
rect 230 1818 234 1822
rect 398 1818 402 1822
rect 782 1818 786 1822
rect 902 1818 906 1822
rect 990 1818 994 1822
rect 1446 1818 1450 1822
rect 1710 1818 1714 1822
rect 1838 1818 1842 1822
rect 2502 1818 2506 1822
rect 2558 1818 2562 1822
rect 2598 1818 2602 1822
rect 3126 1818 3130 1822
rect 3318 1818 3322 1822
rect 3510 1818 3514 1822
rect 3574 1818 3578 1822
rect 3646 1818 3650 1822
rect 3694 1818 3698 1822
rect 3710 1818 3714 1822
rect 3742 1818 3746 1822
rect 346 1803 350 1807
rect 353 1803 357 1807
rect 1362 1803 1366 1807
rect 1369 1803 1373 1807
rect 2386 1803 2390 1807
rect 2393 1803 2397 1807
rect 3410 1803 3414 1807
rect 3417 1803 3421 1807
rect 182 1788 186 1792
rect 454 1788 458 1792
rect 630 1788 634 1792
rect 806 1788 810 1792
rect 870 1788 874 1792
rect 1078 1788 1082 1792
rect 1222 1788 1226 1792
rect 1278 1788 1282 1792
rect 1422 1788 1426 1792
rect 1526 1788 1530 1792
rect 1598 1788 1602 1792
rect 2102 1788 2106 1792
rect 2118 1788 2122 1792
rect 2414 1788 2418 1792
rect 3070 1788 3074 1792
rect 3198 1788 3202 1792
rect 3278 1788 3282 1792
rect 3438 1788 3442 1792
rect 566 1778 570 1782
rect 3166 1778 3170 1782
rect 3558 1778 3562 1782
rect 318 1768 322 1772
rect 438 1768 442 1772
rect 574 1768 578 1772
rect 638 1768 642 1772
rect 814 1768 818 1772
rect 990 1768 994 1772
rect 1566 1768 1570 1772
rect 1926 1768 1930 1772
rect 2262 1768 2266 1772
rect 2694 1768 2698 1772
rect 2878 1768 2882 1772
rect 3174 1768 3178 1772
rect 3478 1768 3482 1772
rect 3550 1768 3554 1772
rect 3582 1768 3586 1772
rect 3614 1768 3618 1772
rect 3662 1768 3666 1772
rect 3678 1768 3682 1772
rect 3710 1768 3714 1772
rect 3758 1768 3762 1772
rect 182 1758 186 1762
rect 326 1758 330 1762
rect 470 1758 474 1762
rect 518 1758 522 1762
rect 550 1758 554 1762
rect 558 1758 562 1762
rect 622 1758 626 1762
rect 654 1758 658 1762
rect 798 1758 802 1762
rect 1006 1758 1010 1762
rect 1222 1758 1226 1762
rect 1246 1758 1250 1762
rect 1422 1758 1426 1762
rect 1478 1758 1482 1762
rect 1502 1758 1506 1762
rect 1550 1758 1554 1762
rect 1582 1758 1586 1762
rect 1622 1758 1626 1762
rect 1638 1758 1642 1762
rect 1782 1758 1786 1762
rect 1814 1758 1818 1762
rect 1894 1758 1898 1762
rect 1998 1758 2002 1762
rect 2070 1758 2074 1762
rect 2414 1758 2418 1762
rect 2454 1758 2458 1762
rect 2470 1758 2474 1762
rect 2486 1758 2490 1762
rect 2518 1758 2522 1762
rect 2550 1758 2554 1762
rect 2582 1758 2586 1762
rect 2614 1758 2618 1762
rect 2678 1758 2682 1762
rect 2710 1758 2714 1762
rect 2766 1758 2770 1762
rect 182 1748 186 1752
rect 294 1748 298 1752
rect 310 1748 314 1752
rect 334 1748 338 1752
rect 358 1748 362 1752
rect 454 1748 458 1752
rect 470 1748 474 1752
rect 502 1748 506 1752
rect 534 1748 538 1752
rect 550 1748 554 1752
rect 566 1748 570 1752
rect 590 1748 594 1752
rect 630 1748 634 1752
rect 654 1748 658 1752
rect 670 1748 674 1752
rect 694 1748 698 1752
rect 766 1748 770 1752
rect 790 1748 794 1752
rect 806 1748 810 1752
rect 838 1748 842 1752
rect 846 1748 850 1752
rect 854 1748 858 1752
rect 886 1748 890 1752
rect 918 1748 922 1752
rect 934 1748 938 1752
rect 950 1748 954 1752
rect 974 1748 978 1752
rect 998 1748 1002 1752
rect 1022 1748 1026 1752
rect 1038 1748 1042 1752
rect 1222 1748 1226 1752
rect 1374 1748 1378 1752
rect 1526 1748 1530 1752
rect 1574 1748 1578 1752
rect 1598 1748 1602 1752
rect 1614 1748 1618 1752
rect 1742 1748 1746 1752
rect 1750 1748 1754 1752
rect 1798 1748 1802 1752
rect 1830 1748 1834 1752
rect 1846 1748 1850 1752
rect 1926 1748 1930 1752
rect 1974 1748 1978 1752
rect 2006 1748 2010 1752
rect 2086 1748 2090 1752
rect 2118 1748 2122 1752
rect 2134 1748 2138 1752
rect 2158 1748 2162 1752
rect 2222 1748 2226 1752
rect 2254 1748 2258 1752
rect 2310 1748 2314 1752
rect 2414 1748 2418 1752
rect 2470 1748 2474 1752
rect 2486 1748 2490 1752
rect 2502 1748 2506 1752
rect 2534 1748 2538 1752
rect 2566 1748 2570 1752
rect 2582 1748 2586 1752
rect 2598 1748 2602 1752
rect 2630 1748 2634 1752
rect 2638 1748 2642 1752
rect 2670 1748 2674 1752
rect 2694 1748 2698 1752
rect 2726 1748 2730 1752
rect 2750 1748 2754 1752
rect 2790 1748 2794 1752
rect 2806 1758 2810 1762
rect 2846 1758 2850 1762
rect 2950 1758 2954 1762
rect 3150 1758 3154 1762
rect 3190 1758 3194 1762
rect 3254 1758 3258 1762
rect 3366 1758 3370 1762
rect 3406 1758 3410 1762
rect 3534 1758 3538 1762
rect 3566 1758 3570 1762
rect 3598 1758 3602 1762
rect 3630 1758 3634 1762
rect 3638 1758 3642 1762
rect 3694 1758 3698 1762
rect 3742 1758 3746 1762
rect 3774 1758 3778 1762
rect 2822 1748 2826 1752
rect 2862 1748 2866 1752
rect 2878 1748 2882 1752
rect 2942 1748 2946 1752
rect 2974 1748 2978 1752
rect 2990 1748 2994 1752
rect 3086 1748 3090 1752
rect 3118 1748 3122 1752
rect 3134 1748 3138 1752
rect 3166 1748 3170 1752
rect 3214 1748 3218 1752
rect 3230 1748 3234 1752
rect 3294 1748 3298 1752
rect 3342 1748 3346 1752
rect 3454 1748 3458 1752
rect 3478 1748 3482 1752
rect 3502 1748 3506 1752
rect 3518 1748 3522 1752
rect 3526 1748 3530 1752
rect 3558 1748 3562 1752
rect 3590 1748 3594 1752
rect 3614 1748 3618 1752
rect 3646 1748 3650 1752
rect 3686 1748 3690 1752
rect 3718 1748 3722 1752
rect 3766 1748 3770 1752
rect 6 1738 10 1742
rect 134 1738 138 1742
rect 270 1738 274 1742
rect 414 1738 418 1742
rect 430 1738 434 1742
rect 446 1738 450 1742
rect 486 1738 490 1742
rect 494 1738 498 1742
rect 510 1738 514 1742
rect 526 1738 530 1742
rect 678 1738 682 1742
rect 686 1738 690 1742
rect 750 1738 754 1742
rect 758 1738 762 1742
rect 790 1738 794 1742
rect 830 1738 834 1742
rect 886 1738 890 1742
rect 910 1738 914 1742
rect 926 1738 930 1742
rect 942 1738 946 1742
rect 998 1738 1002 1742
rect 1030 1738 1034 1742
rect 1062 1738 1066 1742
rect 1174 1738 1178 1742
rect 1262 1738 1266 1742
rect 1374 1738 1378 1742
rect 1454 1738 1458 1742
rect 1486 1738 1490 1742
rect 1518 1738 1522 1742
rect 1574 1738 1578 1742
rect 1606 1738 1610 1742
rect 1614 1738 1618 1742
rect 1646 1738 1650 1742
rect 1710 1738 1714 1742
rect 1726 1738 1730 1742
rect 1758 1738 1762 1742
rect 1806 1738 1810 1742
rect 1838 1738 1842 1742
rect 1854 1738 1858 1742
rect 1910 1738 1914 1742
rect 1918 1738 1922 1742
rect 1966 1738 1970 1742
rect 1982 1738 1986 1742
rect 2006 1738 2010 1742
rect 2014 1738 2018 1742
rect 2030 1738 2034 1742
rect 2062 1738 2066 1742
rect 2094 1738 2098 1742
rect 2110 1738 2114 1742
rect 2198 1738 2202 1742
rect 2246 1738 2250 1742
rect 2366 1738 2370 1742
rect 2478 1738 2482 1742
rect 2510 1738 2514 1742
rect 2542 1738 2546 1742
rect 2574 1738 2578 1742
rect 2606 1738 2610 1742
rect 2638 1738 2642 1742
rect 2662 1738 2666 1742
rect 2702 1738 2706 1742
rect 2734 1738 2738 1742
rect 2742 1738 2746 1742
rect 2774 1738 2778 1742
rect 2830 1738 2834 1742
rect 2870 1738 2874 1742
rect 2934 1738 2938 1742
rect 2966 1738 2970 1742
rect 3030 1738 3034 1742
rect 3094 1738 3098 1742
rect 3110 1738 3114 1742
rect 3126 1738 3130 1742
rect 3206 1738 3210 1742
rect 3222 1738 3226 1742
rect 3238 1738 3242 1742
rect 3270 1738 3274 1742
rect 3302 1738 3306 1742
rect 3334 1738 3338 1742
rect 3350 1738 3354 1742
rect 3382 1738 3386 1742
rect 3390 1738 3394 1742
rect 3734 1738 3738 1742
rect 118 1728 122 1732
rect 278 1728 282 1732
rect 334 1728 338 1732
rect 350 1728 354 1732
rect 422 1728 426 1732
rect 766 1728 770 1732
rect 902 1728 906 1732
rect 990 1728 994 1732
rect 1158 1728 1162 1732
rect 1358 1728 1362 1732
rect 1542 1728 1546 1732
rect 1774 1728 1778 1732
rect 1782 1728 1786 1732
rect 1870 1728 1874 1732
rect 1950 1728 1954 1732
rect 2030 1728 2034 1732
rect 2062 1728 2066 1732
rect 2142 1728 2146 1732
rect 2206 1728 2210 1732
rect 2350 1728 2354 1732
rect 2646 1728 2650 1732
rect 2918 1728 2922 1732
rect 2974 1728 2978 1732
rect 3006 1728 3010 1732
rect 3078 1728 3082 1732
rect 3286 1728 3290 1732
rect 3318 1728 3322 1732
rect 3462 1728 3466 1732
rect 3486 1728 3490 1732
rect 3590 1728 3594 1732
rect 214 1718 218 1722
rect 382 1718 386 1722
rect 606 1718 610 1722
rect 710 1718 714 1722
rect 742 1718 746 1722
rect 1254 1718 1258 1722
rect 1470 1718 1474 1722
rect 1494 1718 1498 1722
rect 1502 1718 1506 1722
rect 1766 1718 1770 1722
rect 1814 1718 1818 1722
rect 1862 1718 1866 1722
rect 1902 1718 1906 1722
rect 2054 1718 2058 1722
rect 2102 1718 2106 1722
rect 2190 1718 2194 1722
rect 2238 1718 2242 1722
rect 2518 1718 2522 1722
rect 2550 1718 2554 1722
rect 2614 1718 2618 1722
rect 2710 1718 2714 1722
rect 3054 1718 3058 1722
rect 3102 1718 3106 1722
rect 3278 1718 3282 1722
rect 3422 1718 3426 1722
rect 3670 1718 3674 1722
rect 3718 1718 3722 1722
rect 3750 1718 3754 1722
rect 850 1703 854 1707
rect 857 1703 861 1707
rect 1882 1703 1886 1707
rect 1889 1703 1893 1707
rect 2906 1703 2910 1707
rect 2913 1703 2917 1707
rect 406 1688 410 1692
rect 582 1688 586 1692
rect 678 1688 682 1692
rect 742 1688 746 1692
rect 822 1688 826 1692
rect 878 1688 882 1692
rect 926 1688 930 1692
rect 950 1688 954 1692
rect 1014 1688 1018 1692
rect 1094 1688 1098 1692
rect 1206 1688 1210 1692
rect 1246 1688 1250 1692
rect 1318 1688 1322 1692
rect 1526 1688 1530 1692
rect 1542 1688 1546 1692
rect 1750 1688 1754 1692
rect 1790 1688 1794 1692
rect 1838 1688 1842 1692
rect 1934 1688 1938 1692
rect 2022 1688 2026 1692
rect 2102 1688 2106 1692
rect 2134 1688 2138 1692
rect 2150 1688 2154 1692
rect 2374 1688 2378 1692
rect 2558 1688 2562 1692
rect 2790 1688 2794 1692
rect 2926 1688 2930 1692
rect 2974 1688 2978 1692
rect 3022 1688 3026 1692
rect 3046 1688 3050 1692
rect 3078 1688 3082 1692
rect 3126 1688 3130 1692
rect 3150 1688 3154 1692
rect 3222 1688 3226 1692
rect 3254 1688 3258 1692
rect 3334 1688 3338 1692
rect 3350 1688 3354 1692
rect 3486 1688 3490 1692
rect 3542 1688 3546 1692
rect 3742 1688 3746 1692
rect 94 1678 98 1682
rect 262 1678 266 1682
rect 366 1678 370 1682
rect 390 1678 394 1682
rect 486 1678 490 1682
rect 942 1678 946 1682
rect 966 1678 970 1682
rect 1006 1678 1010 1682
rect 1054 1678 1058 1682
rect 1070 1678 1074 1682
rect 1254 1678 1258 1682
rect 1374 1678 1378 1682
rect 1486 1678 1490 1682
rect 1518 1678 1522 1682
rect 1638 1678 1642 1682
rect 1822 1678 1826 1682
rect 1918 1678 1922 1682
rect 1942 1678 1946 1682
rect 2030 1678 2034 1682
rect 2062 1678 2066 1682
rect 2078 1678 2082 1682
rect 2230 1678 2234 1682
rect 2318 1678 2322 1682
rect 2358 1678 2362 1682
rect 2454 1678 2458 1682
rect 2598 1678 2602 1682
rect 2654 1678 2658 1682
rect 2678 1678 2682 1682
rect 2782 1678 2786 1682
rect 2814 1678 2818 1682
rect 2846 1678 2850 1682
rect 2886 1678 2890 1682
rect 2982 1678 2986 1682
rect 3006 1678 3010 1682
rect 3142 1678 3146 1682
rect 3214 1678 3218 1682
rect 3270 1678 3274 1682
rect 3286 1678 3290 1682
rect 3342 1678 3346 1682
rect 3374 1678 3378 1682
rect 3398 1678 3402 1682
rect 3430 1678 3434 1682
rect 3494 1678 3498 1682
rect 3550 1678 3554 1682
rect 3574 1678 3578 1682
rect 3630 1678 3634 1682
rect 3654 1678 3658 1682
rect 110 1668 114 1672
rect 246 1668 250 1672
rect 302 1668 306 1672
rect 502 1668 506 1672
rect 590 1668 594 1672
rect 598 1668 602 1672
rect 614 1668 618 1672
rect 662 1668 666 1672
rect 686 1668 690 1672
rect 718 1668 722 1672
rect 750 1668 754 1672
rect 766 1668 770 1672
rect 782 1668 786 1672
rect 158 1658 162 1662
rect 206 1658 210 1662
rect 366 1658 370 1662
rect 446 1658 450 1662
rect 574 1658 578 1662
rect 606 1658 610 1662
rect 638 1658 642 1662
rect 710 1658 714 1662
rect 726 1658 730 1662
rect 758 1658 762 1662
rect 774 1658 778 1662
rect 806 1668 810 1672
rect 846 1668 850 1672
rect 902 1668 906 1672
rect 934 1668 938 1672
rect 1030 1668 1034 1672
rect 1110 1668 1114 1672
rect 1118 1668 1122 1672
rect 1174 1668 1178 1672
rect 1182 1668 1186 1672
rect 1206 1668 1210 1672
rect 1238 1668 1242 1672
rect 1262 1668 1266 1672
rect 1310 1668 1314 1672
rect 1342 1668 1346 1672
rect 1358 1668 1362 1672
rect 1454 1668 1458 1672
rect 1462 1668 1466 1672
rect 1550 1668 1554 1672
rect 1622 1668 1626 1672
rect 1726 1668 1730 1672
rect 1734 1668 1738 1672
rect 1758 1668 1762 1672
rect 1782 1668 1786 1672
rect 1846 1668 1850 1672
rect 1902 1668 1906 1672
rect 1926 1668 1930 1672
rect 1982 1668 1986 1672
rect 1998 1668 2002 1672
rect 2046 1668 2050 1672
rect 2094 1668 2098 1672
rect 2110 1668 2114 1672
rect 2126 1668 2130 1672
rect 2246 1668 2250 1672
rect 2326 1668 2330 1672
rect 2470 1668 2474 1672
rect 2542 1668 2546 1672
rect 2550 1668 2554 1672
rect 2566 1668 2570 1672
rect 2582 1668 2586 1672
rect 2598 1668 2602 1672
rect 2630 1668 2634 1672
rect 2670 1668 2674 1672
rect 2710 1668 2714 1672
rect 2718 1668 2722 1672
rect 2766 1668 2770 1672
rect 2798 1668 2802 1672
rect 2838 1668 2842 1672
rect 2870 1668 2874 1672
rect 2918 1668 2922 1672
rect 2966 1668 2970 1672
rect 3070 1668 3074 1672
rect 3086 1668 3090 1672
rect 3110 1668 3114 1672
rect 3134 1668 3138 1672
rect 3158 1668 3162 1672
rect 3174 1668 3178 1672
rect 3230 1668 3234 1672
rect 3262 1668 3266 1672
rect 3318 1668 3322 1672
rect 3358 1668 3362 1672
rect 3438 1668 3442 1672
rect 3566 1668 3570 1672
rect 3598 1668 3602 1672
rect 3614 1668 3618 1672
rect 3646 1668 3650 1672
rect 3678 1668 3682 1672
rect 798 1658 802 1662
rect 838 1658 842 1662
rect 894 1658 898 1662
rect 910 1658 914 1662
rect 926 1658 930 1662
rect 966 1658 970 1662
rect 982 1658 986 1662
rect 990 1658 994 1662
rect 1038 1658 1042 1662
rect 1086 1658 1090 1662
rect 1230 1658 1234 1662
rect 1270 1658 1274 1662
rect 1334 1658 1338 1662
rect 1350 1658 1354 1662
rect 1366 1658 1370 1662
rect 1382 1658 1386 1662
rect 1414 1658 1418 1662
rect 1502 1658 1506 1662
rect 1574 1658 1578 1662
rect 1766 1658 1770 1662
rect 1774 1658 1778 1662
rect 1806 1658 1810 1662
rect 1854 1658 1858 1662
rect 1870 1658 1874 1662
rect 1894 1658 1898 1662
rect 1910 1658 1914 1662
rect 1958 1658 1962 1662
rect 1990 1658 1994 1662
rect 2006 1658 2010 1662
rect 2054 1658 2058 1662
rect 2062 1658 2066 1662
rect 2078 1658 2082 1662
rect 2118 1658 2122 1662
rect 2246 1658 2250 1662
rect 2294 1658 2298 1662
rect 2414 1658 2418 1662
rect 2510 1658 2514 1662
rect 2526 1658 2530 1662
rect 2574 1658 2578 1662
rect 2622 1658 2626 1662
rect 2638 1658 2642 1662
rect 2702 1658 2706 1662
rect 2726 1658 2730 1662
rect 2774 1658 2778 1662
rect 2814 1658 2818 1662
rect 2830 1658 2834 1662
rect 2870 1658 2874 1662
rect 2910 1658 2914 1662
rect 2958 1658 2962 1662
rect 2982 1658 2986 1662
rect 2990 1658 2994 1662
rect 3038 1658 3042 1662
rect 3166 1658 3170 1662
rect 3238 1658 3242 1662
rect 3286 1658 3290 1662
rect 3310 1658 3314 1662
rect 3366 1658 3370 1662
rect 3390 1658 3394 1662
rect 3414 1658 3418 1662
rect 3454 1658 3458 1662
rect 3470 1658 3474 1662
rect 3518 1658 3522 1662
rect 3526 1658 3530 1662
rect 3566 1658 3570 1662
rect 3590 1658 3594 1662
rect 3598 1658 3602 1662
rect 3646 1658 3650 1662
rect 3654 1658 3658 1662
rect 3670 1658 3674 1662
rect 3686 1658 3690 1662
rect 3694 1658 3698 1662
rect 3726 1658 3730 1662
rect 3758 1658 3762 1662
rect 142 1650 146 1654
rect 214 1650 218 1654
rect 534 1650 538 1654
rect 630 1648 634 1652
rect 742 1648 746 1652
rect 822 1648 826 1652
rect 1142 1648 1146 1652
rect 1158 1648 1162 1652
rect 1198 1648 1202 1652
rect 1286 1648 1290 1652
rect 1398 1648 1402 1652
rect 1430 1648 1434 1652
rect 1478 1648 1482 1652
rect 1486 1648 1490 1652
rect 1590 1650 1594 1654
rect 1886 1648 1890 1652
rect 2294 1648 2298 1652
rect 2502 1650 2506 1654
rect 2686 1648 2690 1652
rect 2742 1648 2746 1652
rect 2814 1648 2818 1652
rect 2942 1648 2946 1652
rect 3046 1648 3050 1652
rect 3086 1648 3090 1652
rect 3094 1648 3098 1652
rect 3118 1648 3122 1652
rect 3246 1648 3250 1652
rect 3334 1648 3338 1652
rect 3486 1648 3490 1652
rect 3542 1648 3546 1652
rect 3622 1648 3626 1652
rect 3702 1648 3706 1652
rect 3734 1648 3738 1652
rect 3766 1648 3770 1652
rect 646 1638 650 1642
rect 678 1638 682 1642
rect 1190 1638 1194 1642
rect 1214 1638 1218 1642
rect 1854 1638 1858 1642
rect 3182 1638 3186 1642
rect 3390 1638 3394 1642
rect 3590 1638 3594 1642
rect 3718 1638 3722 1642
rect 3750 1638 3754 1642
rect 342 1628 346 1632
rect 534 1627 538 1631
rect 1590 1627 1594 1631
rect 2502 1627 2506 1631
rect 3726 1628 3730 1632
rect 14 1618 18 1622
rect 142 1618 146 1622
rect 214 1618 218 1622
rect 670 1618 674 1622
rect 982 1618 986 1622
rect 1166 1618 1170 1622
rect 1966 1618 1970 1622
rect 2294 1618 2298 1622
rect 2702 1618 2706 1622
rect 2750 1618 2754 1622
rect 3286 1618 3290 1622
rect 3310 1618 3314 1622
rect 346 1603 350 1607
rect 353 1603 357 1607
rect 1362 1603 1366 1607
rect 1369 1603 1373 1607
rect 2386 1603 2390 1607
rect 2393 1603 2397 1607
rect 3410 1603 3414 1607
rect 3417 1603 3421 1607
rect 6 1588 10 1592
rect 142 1588 146 1592
rect 454 1588 458 1592
rect 510 1588 514 1592
rect 694 1588 698 1592
rect 758 1588 762 1592
rect 830 1588 834 1592
rect 910 1588 914 1592
rect 942 1588 946 1592
rect 966 1588 970 1592
rect 1006 1588 1010 1592
rect 1158 1588 1162 1592
rect 1230 1588 1234 1592
rect 1374 1588 1378 1592
rect 1422 1588 1426 1592
rect 1494 1588 1498 1592
rect 1518 1588 1522 1592
rect 1574 1588 1578 1592
rect 1598 1588 1602 1592
rect 1630 1588 1634 1592
rect 1774 1588 1778 1592
rect 1942 1588 1946 1592
rect 2118 1588 2122 1592
rect 2262 1588 2266 1592
rect 2286 1588 2290 1592
rect 2358 1588 2362 1592
rect 2502 1588 2506 1592
rect 2670 1588 2674 1592
rect 2686 1588 2690 1592
rect 2830 1588 2834 1592
rect 3174 1588 3178 1592
rect 3198 1588 3202 1592
rect 3534 1588 3538 1592
rect 3670 1588 3674 1592
rect 470 1578 474 1582
rect 1198 1578 1202 1582
rect 2070 1579 2074 1583
rect 30 1568 34 1572
rect 566 1568 570 1572
rect 670 1568 674 1572
rect 702 1568 706 1572
rect 1206 1568 1210 1572
rect 1430 1568 1434 1572
rect 1526 1568 1530 1572
rect 2894 1568 2898 1572
rect 3702 1568 3706 1572
rect 142 1558 146 1562
rect 302 1558 306 1562
rect 326 1558 330 1562
rect 382 1558 386 1562
rect 390 1558 394 1562
rect 486 1558 490 1562
rect 550 1558 554 1562
rect 558 1558 562 1562
rect 582 1558 586 1562
rect 590 1558 594 1562
rect 686 1558 690 1562
rect 750 1558 754 1562
rect 998 1558 1002 1562
rect 1086 1558 1090 1562
rect 1110 1558 1114 1562
rect 1134 1558 1138 1562
rect 1166 1558 1170 1562
rect 1190 1558 1194 1562
rect 1374 1558 1378 1562
rect 1414 1558 1418 1562
rect 1470 1558 1474 1562
rect 22 1548 26 1552
rect 46 1548 50 1552
rect 158 1548 162 1552
rect 438 1548 442 1552
rect 494 1548 498 1552
rect 518 1548 522 1552
rect 574 1548 578 1552
rect 590 1548 594 1552
rect 606 1548 610 1552
rect 622 1548 626 1552
rect 654 1548 658 1552
rect 694 1548 698 1552
rect 718 1548 722 1552
rect 742 1548 746 1552
rect 814 1548 818 1552
rect 862 1548 866 1552
rect 894 1548 898 1552
rect 926 1548 930 1552
rect 958 1548 962 1552
rect 982 1548 986 1552
rect 1046 1548 1050 1552
rect 1054 1548 1058 1552
rect 1206 1548 1210 1552
rect 1270 1548 1274 1552
rect 1430 1548 1434 1552
rect 1454 1548 1458 1552
rect 1510 1558 1514 1562
rect 1774 1558 1778 1562
rect 2070 1556 2074 1560
rect 2262 1558 2266 1562
rect 2502 1558 2506 1562
rect 2582 1558 2586 1562
rect 2622 1558 2626 1562
rect 2654 1558 2658 1562
rect 2830 1558 2834 1562
rect 2854 1558 2858 1562
rect 2910 1558 2914 1562
rect 2998 1558 3002 1562
rect 3014 1558 3018 1562
rect 3110 1558 3114 1562
rect 3166 1558 3170 1562
rect 3190 1558 3194 1562
rect 3214 1558 3218 1562
rect 3494 1558 3498 1562
rect 3550 1558 3554 1562
rect 3590 1558 3594 1562
rect 3622 1558 3626 1562
rect 3718 1558 3722 1562
rect 3734 1558 3738 1562
rect 1494 1548 1498 1552
rect 1526 1548 1530 1552
rect 1614 1548 1618 1552
rect 1766 1548 1770 1552
rect 1814 1548 1818 1552
rect 1878 1548 1882 1552
rect 1886 1548 1890 1552
rect 118 1538 122 1542
rect 190 1538 194 1542
rect 318 1538 322 1542
rect 342 1538 346 1542
rect 366 1538 370 1542
rect 406 1538 410 1542
rect 430 1538 434 1542
rect 446 1538 450 1542
rect 462 1538 466 1542
rect 526 1538 530 1542
rect 2086 1548 2090 1552
rect 2246 1548 2250 1552
rect 2302 1548 2306 1552
rect 2502 1548 2506 1552
rect 2526 1548 2530 1552
rect 2550 1548 2554 1552
rect 2614 1548 2618 1552
rect 2638 1548 2642 1552
rect 2726 1548 2730 1552
rect 2870 1548 2874 1552
rect 2878 1548 2882 1552
rect 2934 1548 2938 1552
rect 2990 1548 2994 1552
rect 3022 1548 3026 1552
rect 3030 1548 3034 1552
rect 3046 1548 3050 1552
rect 3054 1548 3058 1552
rect 3078 1548 3082 1552
rect 3126 1548 3130 1552
rect 3142 1548 3146 1552
rect 3254 1548 3258 1552
rect 3278 1548 3282 1552
rect 3286 1548 3290 1552
rect 3318 1548 3322 1552
rect 3350 1548 3354 1552
rect 3358 1548 3362 1552
rect 3390 1548 3394 1552
rect 3398 1548 3402 1552
rect 3430 1548 3434 1552
rect 3454 1548 3458 1552
rect 3486 1548 3490 1552
rect 3510 1548 3514 1552
rect 3542 1548 3546 1552
rect 3582 1548 3586 1552
rect 3606 1548 3610 1552
rect 3638 1548 3642 1552
rect 3686 1548 3690 1552
rect 3710 1548 3714 1552
rect 3750 1548 3754 1552
rect 614 1538 618 1542
rect 638 1538 642 1542
rect 718 1538 722 1542
rect 790 1538 794 1542
rect 958 1538 962 1542
rect 990 1538 994 1542
rect 1014 1538 1018 1542
rect 1102 1538 1106 1542
rect 1126 1538 1130 1542
rect 1150 1538 1154 1542
rect 1326 1538 1330 1542
rect 1446 1538 1450 1542
rect 1502 1538 1506 1542
rect 1558 1538 1562 1542
rect 1726 1538 1730 1542
rect 1838 1538 1842 1542
rect 1870 1538 1874 1542
rect 1982 1538 1986 1542
rect 2038 1538 2042 1542
rect 2214 1538 2218 1542
rect 2294 1538 2298 1542
rect 2326 1538 2330 1542
rect 2454 1538 2458 1542
rect 2566 1538 2570 1542
rect 2606 1538 2610 1542
rect 2646 1538 2650 1542
rect 2662 1538 2666 1542
rect 2782 1538 2786 1542
rect 2878 1538 2882 1542
rect 2886 1538 2890 1542
rect 2982 1538 2986 1542
rect 3086 1538 3090 1542
rect 3134 1538 3138 1542
rect 3182 1538 3186 1542
rect 3206 1538 3210 1542
rect 3230 1538 3234 1542
rect 3294 1538 3298 1542
rect 3310 1538 3314 1542
rect 3342 1538 3346 1542
rect 3366 1538 3370 1542
rect 3374 1538 3378 1542
rect 3382 1538 3386 1542
rect 3406 1538 3410 1542
rect 3422 1538 3426 1542
rect 3462 1538 3466 1542
rect 3470 1538 3474 1542
rect 3486 1538 3490 1542
rect 3526 1538 3530 1542
rect 3614 1538 3618 1542
rect 206 1528 210 1532
rect 286 1528 290 1532
rect 414 1528 418 1532
rect 750 1528 754 1532
rect 766 1528 770 1532
rect 806 1528 810 1532
rect 830 1528 834 1532
rect 1030 1528 1034 1532
rect 1166 1528 1170 1532
rect 1182 1528 1186 1532
rect 1310 1528 1314 1532
rect 1542 1528 1546 1532
rect 1566 1528 1570 1532
rect 1582 1528 1586 1532
rect 1710 1528 1714 1532
rect 1798 1528 1802 1532
rect 1830 1528 1834 1532
rect 1854 1528 1858 1532
rect 1918 1528 1922 1532
rect 2022 1528 2026 1532
rect 2198 1528 2202 1532
rect 2438 1528 2442 1532
rect 2542 1528 2546 1532
rect 2766 1528 2770 1532
rect 2854 1528 2858 1532
rect 2966 1528 2970 1532
rect 3046 1528 3050 1532
rect 3070 1528 3074 1532
rect 3158 1528 3162 1532
rect 3238 1528 3242 1532
rect 3262 1528 3266 1532
rect 3326 1528 3330 1532
rect 3526 1528 3530 1532
rect 3542 1528 3546 1532
rect 3622 1528 3626 1532
rect 3638 1528 3642 1532
rect 3654 1528 3658 1532
rect 62 1518 66 1522
rect 310 1518 314 1522
rect 326 1518 330 1522
rect 382 1518 386 1522
rect 390 1518 394 1522
rect 422 1518 426 1522
rect 550 1518 554 1522
rect 798 1518 802 1522
rect 878 1518 882 1522
rect 910 1518 914 1522
rect 942 1518 946 1522
rect 1070 1518 1074 1522
rect 1094 1518 1098 1522
rect 1118 1518 1122 1522
rect 1142 1518 1146 1522
rect 2950 1518 2954 1522
rect 2974 1518 2978 1522
rect 3094 1518 3098 1522
rect 3150 1518 3154 1522
rect 3214 1518 3218 1522
rect 3246 1518 3250 1522
rect 3270 1518 3274 1522
rect 3310 1518 3314 1522
rect 3334 1518 3338 1522
rect 3422 1518 3426 1522
rect 3494 1518 3498 1522
rect 3574 1518 3578 1522
rect 3590 1518 3594 1522
rect 3670 1518 3674 1522
rect 3702 1518 3706 1522
rect 850 1503 854 1507
rect 857 1503 861 1507
rect 1882 1503 1886 1507
rect 1889 1503 1893 1507
rect 2906 1503 2910 1507
rect 2913 1503 2917 1507
rect 510 1488 514 1492
rect 542 1488 546 1492
rect 710 1488 714 1492
rect 726 1488 730 1492
rect 766 1488 770 1492
rect 998 1488 1002 1492
rect 1022 1488 1026 1492
rect 1102 1488 1106 1492
rect 1142 1488 1146 1492
rect 1286 1488 1290 1492
rect 1326 1488 1330 1492
rect 1366 1488 1370 1492
rect 1782 1488 1786 1492
rect 1830 1488 1834 1492
rect 1878 1488 1882 1492
rect 1958 1488 1962 1492
rect 2150 1488 2154 1492
rect 2366 1488 2370 1492
rect 2526 1488 2530 1492
rect 2582 1488 2586 1492
rect 2606 1488 2610 1492
rect 2886 1488 2890 1492
rect 3182 1488 3186 1492
rect 3614 1488 3618 1492
rect 3694 1488 3698 1492
rect 86 1478 90 1482
rect 262 1478 266 1482
rect 366 1478 370 1482
rect 382 1478 386 1482
rect 454 1478 458 1482
rect 518 1478 522 1482
rect 630 1478 634 1482
rect 1046 1478 1050 1482
rect 1094 1478 1098 1482
rect 1150 1478 1154 1482
rect 1446 1478 1450 1482
rect 1638 1478 1642 1482
rect 1942 1478 1946 1482
rect 2038 1478 2042 1482
rect 2230 1478 2234 1482
rect 2814 1478 2818 1482
rect 2958 1478 2962 1482
rect 3054 1478 3058 1482
rect 3134 1478 3138 1482
rect 3158 1478 3162 1482
rect 3174 1478 3178 1482
rect 3190 1478 3194 1482
rect 3222 1478 3226 1482
rect 3230 1478 3234 1482
rect 3262 1478 3266 1482
rect 3294 1478 3298 1482
rect 3398 1478 3402 1482
rect 3478 1478 3482 1482
rect 3542 1478 3546 1482
rect 3558 1478 3562 1482
rect 3622 1478 3626 1482
rect 3646 1478 3650 1482
rect 3662 1478 3666 1482
rect 70 1468 74 1472
rect 246 1468 250 1472
rect 390 1468 394 1472
rect 422 1468 426 1472
rect 446 1468 450 1472
rect 462 1468 466 1472
rect 478 1468 482 1472
rect 494 1468 498 1472
rect 502 1468 506 1472
rect 534 1468 538 1472
rect 614 1468 618 1472
rect 742 1468 746 1472
rect 838 1468 842 1472
rect 862 1468 866 1472
rect 870 1468 874 1472
rect 934 1468 938 1472
rect 966 1468 970 1472
rect 974 1468 978 1472
rect 1006 1468 1010 1472
rect 1014 1468 1018 1472
rect 1030 1468 1034 1472
rect 1054 1468 1058 1472
rect 1086 1468 1090 1472
rect 1134 1468 1138 1472
rect 1150 1468 1154 1472
rect 1174 1468 1178 1472
rect 1190 1468 1194 1472
rect 1230 1468 1234 1472
rect 1302 1468 1306 1472
rect 1350 1468 1354 1472
rect 1462 1468 1466 1472
rect 1534 1468 1538 1472
rect 1654 1468 1658 1472
rect 1726 1468 1730 1472
rect 1742 1468 1746 1472
rect 1758 1468 1762 1472
rect 1806 1468 1810 1472
rect 1822 1468 1826 1472
rect 1870 1468 1874 1472
rect 1918 1468 1922 1472
rect 2054 1468 2058 1472
rect 2126 1468 2130 1472
rect 2246 1468 2250 1472
rect 2318 1468 2322 1472
rect 2342 1468 2346 1472
rect 2350 1468 2354 1472
rect 2390 1468 2394 1472
rect 2438 1468 2442 1472
rect 2470 1468 2474 1472
rect 2518 1468 2522 1472
rect 2566 1468 2570 1472
rect 2590 1468 2594 1472
rect 2598 1468 2602 1472
rect 2614 1468 2618 1472
rect 126 1458 130 1462
rect 206 1458 210 1462
rect 398 1458 402 1462
rect 470 1458 474 1462
rect 486 1458 490 1462
rect 534 1458 538 1462
rect 574 1458 578 1462
rect 750 1458 754 1462
rect 798 1458 802 1462
rect 814 1458 818 1462
rect 830 1458 834 1462
rect 846 1458 850 1462
rect 918 1458 922 1462
rect 966 1458 970 1462
rect 998 1458 1002 1462
rect 1062 1458 1066 1462
rect 1086 1458 1090 1462
rect 1118 1458 1122 1462
rect 1126 1458 1130 1462
rect 1166 1458 1170 1462
rect 1182 1458 1186 1462
rect 1198 1458 1202 1462
rect 1222 1458 1226 1462
rect 1310 1458 1314 1462
rect 1326 1458 1330 1462
rect 1406 1458 1410 1462
rect 1557 1458 1561 1462
rect 1702 1458 1706 1462
rect 1798 1458 1802 1462
rect 1814 1458 1818 1462
rect 1862 1458 1866 1462
rect 1910 1458 1914 1462
rect 1926 1458 1930 1462
rect 2102 1458 2106 1462
rect 2190 1458 2194 1462
rect 2278 1458 2282 1462
rect 2318 1458 2322 1462
rect 2462 1458 2466 1462
rect 2478 1458 2482 1462
rect 2510 1458 2514 1462
rect 2558 1458 2562 1462
rect 2638 1466 2642 1470
rect 2646 1468 2650 1472
rect 2678 1468 2682 1472
rect 2710 1468 2714 1472
rect 2742 1468 2746 1472
rect 2750 1468 2754 1472
rect 2806 1468 2810 1472
rect 2838 1468 2842 1472
rect 2846 1468 2850 1472
rect 2942 1468 2946 1472
rect 3006 1468 3010 1472
rect 3030 1468 3034 1472
rect 3110 1468 3114 1472
rect 3118 1468 3122 1472
rect 3206 1468 3210 1472
rect 3246 1468 3250 1472
rect 3286 1468 3290 1472
rect 3302 1468 3306 1472
rect 3390 1468 3394 1472
rect 3414 1468 3418 1472
rect 3446 1468 3450 1472
rect 3494 1468 3498 1472
rect 3638 1468 3642 1472
rect 3670 1468 3674 1472
rect 3718 1468 3722 1472
rect 2678 1458 2682 1462
rect 2734 1458 2738 1462
rect 2758 1458 2762 1462
rect 2798 1458 2802 1462
rect 2846 1458 2850 1462
rect 2854 1458 2858 1462
rect 2926 1458 2930 1462
rect 2974 1458 2978 1462
rect 2982 1458 2986 1462
rect 3014 1458 3018 1462
rect 3038 1458 3042 1462
rect 3062 1458 3066 1462
rect 3078 1458 3082 1462
rect 3086 1458 3090 1462
rect 3118 1458 3122 1462
rect 3142 1458 3146 1462
rect 3158 1458 3162 1462
rect 3198 1458 3202 1462
rect 3294 1458 3298 1462
rect 3358 1458 3362 1462
rect 3366 1458 3370 1462
rect 3422 1458 3426 1462
rect 3454 1458 3458 1462
rect 3502 1458 3506 1462
rect 3534 1458 3538 1462
rect 3550 1458 3554 1462
rect 3558 1458 3562 1462
rect 3582 1458 3586 1462
rect 3590 1458 3594 1462
rect 3638 1458 3642 1462
rect 3662 1458 3666 1462
rect 3678 1458 3682 1462
rect 3702 1458 3706 1462
rect 3758 1458 3762 1462
rect 14 1448 18 1452
rect 198 1448 202 1452
rect 398 1448 402 1452
rect 430 1448 434 1452
rect 566 1448 570 1452
rect 806 1448 810 1452
rect 814 1448 818 1452
rect 950 1448 954 1452
rect 1078 1448 1082 1452
rect 1510 1448 1514 1452
rect 1702 1448 1706 1452
rect 1774 1448 1778 1452
rect 1846 1448 1850 1452
rect 1894 1448 1898 1452
rect 1934 1448 1938 1452
rect 2086 1450 2090 1454
rect 2294 1448 2298 1452
rect 2366 1448 2370 1452
rect 2398 1448 2402 1452
rect 2446 1448 2450 1452
rect 2542 1448 2546 1452
rect 2654 1448 2658 1452
rect 2686 1448 2690 1452
rect 2718 1448 2722 1452
rect 2774 1448 2778 1452
rect 2782 1448 2786 1452
rect 2814 1448 2818 1452
rect 2854 1448 2858 1452
rect 2870 1448 2874 1452
rect 3014 1448 3018 1452
rect 3614 1448 3618 1452
rect 3694 1448 3698 1452
rect 726 1438 730 1442
rect 790 1438 794 1442
rect 1030 1438 1034 1442
rect 2494 1438 2498 1442
rect 2670 1438 2674 1442
rect 2798 1438 2802 1442
rect 126 1427 130 1431
rect 854 1428 858 1432
rect 958 1428 962 1432
rect 2358 1428 2362 1432
rect 3742 1428 3746 1432
rect 166 1418 170 1422
rect 198 1418 202 1422
rect 374 1418 378 1422
rect 566 1418 570 1422
rect 734 1418 738 1422
rect 798 1418 802 1422
rect 894 1418 898 1422
rect 1510 1418 1514 1422
rect 1542 1418 1546 1422
rect 1702 1418 1706 1422
rect 1734 1418 1738 1422
rect 1750 1418 1754 1422
rect 2086 1418 2090 1422
rect 2134 1418 2138 1422
rect 2294 1418 2298 1422
rect 2702 1418 2706 1422
rect 2758 1418 2762 1422
rect 2966 1418 2970 1422
rect 3038 1418 3042 1422
rect 3166 1418 3170 1422
rect 3222 1418 3226 1422
rect 3342 1418 3346 1422
rect 3398 1418 3402 1422
rect 3454 1418 3458 1422
rect 346 1403 350 1407
rect 353 1403 357 1407
rect 1362 1403 1366 1407
rect 1369 1403 1373 1407
rect 2386 1403 2390 1407
rect 2393 1403 2397 1407
rect 3410 1403 3414 1407
rect 3417 1403 3421 1407
rect 222 1388 226 1392
rect 254 1388 258 1392
rect 518 1388 522 1392
rect 598 1388 602 1392
rect 654 1388 658 1392
rect 878 1388 882 1392
rect 1166 1388 1170 1392
rect 1198 1388 1202 1392
rect 1358 1388 1362 1392
rect 1566 1388 1570 1392
rect 1710 1388 1714 1392
rect 1790 1388 1794 1392
rect 1822 1388 1826 1392
rect 1870 1388 1874 1392
rect 1910 1388 1914 1392
rect 2054 1388 2058 1392
rect 2230 1388 2234 1392
rect 2606 1388 2610 1392
rect 2750 1388 2754 1392
rect 3326 1388 3330 1392
rect 3470 1388 3474 1392
rect 3542 1388 3546 1392
rect 3718 1388 3722 1392
rect 46 1378 50 1382
rect 350 1379 354 1383
rect 486 1368 490 1372
rect 550 1368 554 1372
rect 574 1368 578 1372
rect 1038 1379 1042 1383
rect 1478 1378 1482 1382
rect 3118 1378 3122 1382
rect 718 1368 722 1372
rect 806 1368 810 1372
rect 1646 1368 1650 1372
rect 1742 1368 1746 1372
rect 2118 1368 2122 1372
rect 2286 1368 2290 1372
rect 2854 1368 2858 1372
rect 3462 1368 3466 1372
rect 3694 1368 3698 1372
rect 3702 1368 3706 1372
rect 3726 1368 3730 1372
rect 222 1358 226 1362
rect 270 1358 274 1362
rect 278 1358 282 1362
rect 350 1356 354 1360
rect 534 1358 538 1362
rect 702 1358 706 1362
rect 734 1358 738 1362
rect 822 1358 826 1362
rect 854 1358 858 1362
rect 942 1358 946 1362
rect 1038 1356 1042 1360
rect 1198 1358 1202 1362
rect 1406 1358 1410 1362
rect 222 1348 226 1352
rect 246 1348 250 1352
rect 334 1348 338 1352
rect 526 1348 530 1352
rect 542 1348 546 1352
rect 582 1348 586 1352
rect 590 1348 594 1352
rect 678 1348 682 1352
rect 718 1348 722 1352
rect 750 1348 754 1352
rect 774 1348 778 1352
rect 814 1348 818 1352
rect 830 1348 834 1352
rect 894 1348 898 1352
rect 918 1348 922 1352
rect 958 1348 962 1352
rect 974 1348 978 1352
rect 998 1348 1002 1352
rect 1126 1348 1130 1352
rect 1206 1348 1210 1352
rect 1446 1358 1450 1362
rect 1494 1358 1498 1362
rect 1550 1358 1554 1362
rect 1430 1348 1434 1352
rect 1438 1348 1442 1352
rect 1462 1348 1466 1352
rect 1502 1348 1506 1352
rect 1510 1348 1514 1352
rect 1526 1348 1530 1352
rect 1566 1348 1570 1352
rect 1606 1358 1610 1362
rect 1622 1348 1626 1352
rect 1646 1348 1650 1352
rect 1670 1358 1674 1362
rect 1774 1358 1778 1362
rect 1806 1358 1810 1362
rect 1838 1358 1842 1362
rect 2054 1358 2058 1362
rect 2094 1358 2098 1362
rect 1686 1348 1690 1352
rect 1710 1348 1714 1352
rect 1726 1348 1730 1352
rect 1766 1348 1770 1352
rect 1790 1348 1794 1352
rect 1854 1348 1858 1352
rect 2046 1348 2050 1352
rect 2134 1358 2138 1362
rect 2166 1358 2170 1362
rect 2182 1348 2186 1352
rect 2198 1348 2202 1352
rect 2222 1348 2226 1352
rect 2254 1348 2258 1352
rect 2294 1358 2298 1362
rect 2326 1358 2330 1362
rect 2358 1358 2362 1362
rect 2430 1358 2434 1362
rect 2374 1348 2378 1352
rect 2398 1348 2402 1352
rect 2470 1358 2474 1362
rect 2502 1358 2506 1362
rect 2534 1358 2538 1362
rect 2566 1358 2570 1362
rect 2750 1358 2754 1362
rect 2774 1358 2778 1362
rect 2806 1358 2810 1362
rect 2838 1358 2842 1362
rect 2902 1358 2906 1362
rect 2974 1358 2978 1362
rect 3006 1358 3010 1362
rect 3142 1358 3146 1362
rect 3254 1358 3258 1362
rect 3302 1358 3306 1362
rect 3390 1358 3394 1362
rect 3454 1358 3458 1362
rect 3558 1358 3562 1362
rect 3646 1358 3650 1362
rect 3710 1358 3714 1362
rect 3742 1358 3746 1362
rect 3774 1358 3778 1362
rect 2518 1348 2522 1352
rect 2550 1348 2554 1352
rect 2590 1348 2594 1352
rect 2646 1348 2650 1352
rect 2734 1348 2738 1352
rect 2790 1348 2794 1352
rect 2806 1348 2810 1352
rect 2838 1348 2842 1352
rect 2854 1348 2858 1352
rect 2870 1348 2874 1352
rect 2934 1348 2938 1352
rect 2966 1348 2970 1352
rect 2990 1348 2994 1352
rect 3022 1348 3026 1352
rect 3062 1348 3066 1352
rect 3070 1348 3074 1352
rect 3102 1348 3106 1352
rect 3174 1348 3178 1352
rect 3182 1348 3186 1352
rect 3206 1348 3210 1352
rect 38 1338 42 1342
rect 174 1338 178 1342
rect 246 1338 250 1342
rect 294 1338 298 1342
rect 382 1338 386 1342
rect 510 1338 514 1342
rect 630 1338 634 1342
rect 670 1338 674 1342
rect 734 1338 738 1342
rect 758 1338 762 1342
rect 766 1338 770 1342
rect 830 1338 834 1342
rect 902 1338 906 1342
rect 918 1338 922 1342
rect 926 1338 930 1342
rect 950 1338 954 1342
rect 982 1338 986 1342
rect 1070 1338 1074 1342
rect 1246 1338 1250 1342
rect 1390 1338 1394 1342
rect 1406 1338 1410 1342
rect 1438 1338 1442 1342
rect 1486 1338 1490 1342
rect 1518 1338 1522 1342
rect 1526 1338 1530 1342
rect 1574 1338 1578 1342
rect 1630 1338 1634 1342
rect 1638 1338 1642 1342
rect 1694 1338 1698 1342
rect 1702 1338 1706 1342
rect 1742 1338 1746 1342
rect 1758 1338 1762 1342
rect 1798 1338 1802 1342
rect 1830 1338 1834 1342
rect 1862 1338 1866 1342
rect 2006 1338 2010 1342
rect 2078 1338 2082 1342
rect 2126 1338 2130 1342
rect 2158 1338 2162 1342
rect 2190 1338 2194 1342
rect 2246 1338 2250 1342
rect 2270 1338 2274 1342
rect 2278 1338 2282 1342
rect 2318 1338 2322 1342
rect 2350 1338 2354 1342
rect 2382 1338 2386 1342
rect 2406 1338 2410 1342
rect 2462 1338 2466 1342
rect 2494 1338 2498 1342
rect 2526 1338 2530 1342
rect 2542 1338 2546 1342
rect 2558 1338 2562 1342
rect 2582 1338 2586 1342
rect 2702 1338 2706 1342
rect 2798 1338 2802 1342
rect 2830 1338 2834 1342
rect 2862 1338 2866 1342
rect 2878 1338 2882 1342
rect 2942 1338 2946 1342
rect 2998 1338 3002 1342
rect 3014 1338 3018 1342
rect 3030 1338 3034 1342
rect 3054 1338 3058 1342
rect 3262 1348 3266 1352
rect 3342 1348 3346 1352
rect 3398 1348 3402 1352
rect 3454 1348 3458 1352
rect 3502 1348 3506 1352
rect 3526 1348 3530 1352
rect 3542 1348 3546 1352
rect 3566 1348 3570 1352
rect 3598 1348 3602 1352
rect 3102 1338 3106 1342
rect 3110 1338 3114 1342
rect 3126 1338 3130 1342
rect 3150 1338 3154 1342
rect 3214 1338 3218 1342
rect 3230 1338 3234 1342
rect 3238 1338 3242 1342
rect 3294 1338 3298 1342
rect 3318 1338 3322 1342
rect 3334 1338 3338 1342
rect 3350 1338 3354 1342
rect 3374 1338 3378 1342
rect 3406 1338 3410 1342
rect 3534 1338 3538 1342
rect 3574 1338 3578 1342
rect 158 1328 162 1332
rect 398 1328 402 1332
rect 502 1328 506 1332
rect 510 1328 514 1332
rect 542 1328 546 1332
rect 566 1328 570 1332
rect 998 1328 1002 1332
rect 1086 1328 1090 1332
rect 1262 1328 1266 1332
rect 1342 1328 1346 1332
rect 1374 1328 1378 1332
rect 3630 1348 3634 1352
rect 3646 1348 3650 1352
rect 3702 1348 3706 1352
rect 3734 1348 3738 1352
rect 3758 1348 3762 1352
rect 3774 1348 3778 1352
rect 3622 1338 3626 1342
rect 3646 1338 3650 1342
rect 3678 1338 3682 1342
rect 3750 1338 3754 1342
rect 1542 1328 1546 1332
rect 1590 1328 1594 1332
rect 1742 1328 1746 1332
rect 1902 1328 1906 1332
rect 1990 1328 1994 1332
rect 2238 1328 2242 1332
rect 2566 1328 2570 1332
rect 2686 1328 2690 1332
rect 2950 1328 2954 1332
rect 3038 1328 3042 1332
rect 3086 1328 3090 1332
rect 3198 1328 3202 1332
rect 3230 1328 3234 1332
rect 3366 1328 3370 1332
rect 3422 1328 3426 1332
rect 3510 1328 3514 1332
rect 3590 1328 3594 1332
rect 3598 1328 3602 1332
rect 3614 1328 3618 1332
rect 30 1318 34 1322
rect 278 1318 282 1322
rect 694 1318 698 1322
rect 790 1318 794 1322
rect 870 1318 874 1322
rect 934 1318 938 1322
rect 974 1318 978 1322
rect 2294 1318 2298 1322
rect 2438 1318 2442 1322
rect 2774 1318 2778 1322
rect 2886 1318 2890 1322
rect 2974 1318 2978 1322
rect 3046 1318 3050 1322
rect 3134 1318 3138 1322
rect 3190 1318 3194 1322
rect 3278 1318 3282 1322
rect 3358 1318 3362 1322
rect 3390 1318 3394 1322
rect 3414 1318 3418 1322
rect 3486 1318 3490 1322
rect 3518 1318 3522 1322
rect 3582 1318 3586 1322
rect 850 1303 854 1307
rect 857 1303 861 1307
rect 1882 1303 1886 1307
rect 1889 1303 1893 1307
rect 2906 1303 2910 1307
rect 2913 1303 2917 1307
rect 14 1288 18 1292
rect 118 1288 122 1292
rect 246 1288 250 1292
rect 302 1288 306 1292
rect 542 1288 546 1292
rect 782 1288 786 1292
rect 966 1288 970 1292
rect 990 1288 994 1292
rect 1006 1288 1010 1292
rect 1062 1288 1066 1292
rect 1382 1288 1386 1292
rect 1446 1288 1450 1292
rect 1542 1288 1546 1292
rect 1718 1288 1722 1292
rect 1734 1288 1738 1292
rect 1758 1288 1762 1292
rect 1790 1288 1794 1292
rect 1838 1288 1842 1292
rect 2038 1288 2042 1292
rect 2070 1288 2074 1292
rect 2254 1288 2258 1292
rect 2358 1288 2362 1292
rect 2478 1288 2482 1292
rect 2534 1288 2538 1292
rect 2558 1288 2562 1292
rect 2646 1288 2650 1292
rect 2822 1288 2826 1292
rect 3086 1288 3090 1292
rect 3294 1288 3298 1292
rect 3310 1288 3314 1292
rect 3462 1288 3466 1292
rect 3550 1288 3554 1292
rect 3574 1288 3578 1292
rect 3606 1288 3610 1292
rect 3646 1288 3650 1292
rect 182 1278 186 1282
rect 382 1278 386 1282
rect 470 1278 474 1282
rect 590 1278 594 1282
rect 686 1278 690 1282
rect 886 1278 890 1282
rect 982 1278 986 1282
rect 1054 1278 1058 1282
rect 1086 1278 1090 1282
rect 1142 1278 1146 1282
rect 1158 1278 1162 1282
rect 1270 1278 1274 1282
rect 1350 1278 1354 1282
rect 1390 1278 1394 1282
rect 1414 1278 1418 1282
rect 1470 1278 1474 1282
rect 1534 1278 1538 1282
rect 1582 1278 1586 1282
rect 1726 1278 1730 1282
rect 1918 1278 1922 1282
rect 38 1268 42 1272
rect 102 1268 106 1272
rect 174 1268 178 1272
rect 270 1268 274 1272
rect 398 1268 402 1272
rect 486 1268 490 1272
rect 502 1268 506 1272
rect 534 1268 538 1272
rect 558 1268 562 1272
rect 582 1268 586 1272
rect 702 1268 706 1272
rect 774 1268 778 1272
rect 870 1268 874 1272
rect 1030 1268 1034 1272
rect 1102 1268 1106 1272
rect 1118 1268 1122 1272
rect 1150 1268 1154 1272
rect 1174 1268 1178 1272
rect 1254 1268 1258 1272
rect 1454 1268 1458 1272
rect 1526 1268 1530 1272
rect 1550 1268 1554 1272
rect 1566 1268 1570 1272
rect 1598 1268 1602 1272
rect 1614 1268 1618 1272
rect 1710 1268 1714 1272
rect 1750 1268 1754 1272
rect 1774 1268 1778 1272
rect 1934 1268 1938 1272
rect 2150 1278 2154 1282
rect 2350 1278 2354 1282
rect 2494 1278 2498 1282
rect 2550 1278 2554 1282
rect 2726 1278 2730 1282
rect 2958 1278 2962 1282
rect 3094 1278 3098 1282
rect 3214 1278 3218 1282
rect 3230 1278 3234 1282
rect 3302 1278 3306 1282
rect 3358 1278 3362 1282
rect 3558 1278 3562 1282
rect 3710 1278 3714 1282
rect 2166 1268 2170 1272
rect 2246 1268 2250 1272
rect 2294 1268 2298 1272
rect 2326 1268 2330 1272
rect 2334 1268 2338 1272
rect 2366 1268 2370 1272
rect 2374 1268 2378 1272
rect 2422 1268 2426 1272
rect 2446 1268 2450 1272
rect 2742 1268 2746 1272
rect 2814 1268 2818 1272
rect 2830 1268 2834 1272
rect 2910 1268 2914 1272
rect 2942 1268 2946 1272
rect 2982 1268 2986 1272
rect 3014 1268 3018 1272
rect 3078 1268 3082 1272
rect 3126 1268 3130 1272
rect 3166 1268 3170 1272
rect 3238 1268 3242 1272
rect 3286 1268 3290 1272
rect 3326 1268 3330 1272
rect 3342 1268 3346 1272
rect 3374 1268 3378 1272
rect 3398 1268 3402 1272
rect 3422 1268 3426 1272
rect 3454 1268 3458 1272
rect 3470 1268 3474 1272
rect 3502 1268 3506 1272
rect 3510 1268 3514 1272
rect 3542 1268 3546 1272
rect 3566 1268 3570 1272
rect 3590 1268 3594 1272
rect 3662 1268 3666 1272
rect 3678 1268 3682 1272
rect 3726 1268 3730 1272
rect 3742 1268 3746 1272
rect 3758 1268 3762 1272
rect 30 1258 34 1262
rect 222 1258 226 1262
rect 230 1258 234 1262
rect 342 1258 346 1262
rect 454 1258 458 1262
rect 494 1258 498 1262
rect 566 1258 570 1262
rect 646 1258 650 1262
rect 750 1258 754 1262
rect 822 1258 826 1262
rect 998 1258 1002 1262
rect 1022 1258 1026 1262
rect 1038 1258 1042 1262
rect 1118 1258 1122 1262
rect 1126 1258 1130 1262
rect 1142 1258 1146 1262
rect 1182 1258 1186 1262
rect 1206 1258 1210 1262
rect 1430 1258 1434 1262
rect 1502 1258 1506 1262
rect 1518 1258 1522 1262
rect 1558 1258 1562 1262
rect 1606 1258 1610 1262
rect 1638 1258 1642 1262
rect 1806 1258 1810 1262
rect 1982 1258 1986 1262
rect 2006 1258 2010 1262
rect 2022 1258 2026 1262
rect 2054 1258 2058 1262
rect 2110 1258 2114 1262
rect 2238 1258 2242 1262
rect 2286 1258 2290 1262
rect 2318 1258 2322 1262
rect 2382 1258 2386 1262
rect 2414 1258 2418 1262
rect 2422 1258 2426 1262
rect 2462 1258 2466 1262
rect 2486 1258 2490 1262
rect 2510 1258 2514 1262
rect 2518 1258 2522 1262
rect 2566 1258 2570 1262
rect 2574 1258 2578 1262
rect 2614 1258 2618 1262
rect 2686 1258 2690 1262
rect 2838 1258 2842 1262
rect 2902 1258 2906 1262
rect 2934 1258 2938 1262
rect 2958 1258 2962 1262
rect 2974 1258 2978 1262
rect 3070 1258 3074 1262
rect 3102 1258 3106 1262
rect 3142 1258 3146 1262
rect 3190 1258 3194 1262
rect 3238 1258 3242 1262
rect 3278 1258 3282 1262
rect 3334 1258 3338 1262
rect 3446 1258 3450 1262
rect 3478 1258 3482 1262
rect 3494 1258 3498 1262
rect 3630 1258 3634 1262
rect 3670 1258 3674 1262
rect 3702 1258 3706 1262
rect 3734 1258 3738 1262
rect 214 1248 218 1252
rect 254 1248 258 1252
rect 446 1248 450 1252
rect 518 1248 522 1252
rect 534 1248 538 1252
rect 734 1250 738 1254
rect 838 1250 842 1254
rect 1006 1248 1010 1252
rect 1222 1250 1226 1254
rect 1406 1248 1410 1252
rect 1502 1248 1506 1252
rect 1734 1248 1738 1252
rect 1758 1248 1762 1252
rect 1982 1248 1986 1252
rect 2198 1250 2202 1254
rect 2270 1248 2274 1252
rect 2302 1248 2306 1252
rect 2398 1248 2402 1252
rect 2638 1248 2642 1252
rect 2774 1250 2778 1254
rect 2854 1248 2858 1252
rect 3006 1248 3010 1252
rect 3054 1248 3058 1252
rect 3158 1248 3162 1252
rect 3190 1248 3194 1252
rect 3310 1248 3314 1252
rect 3406 1248 3410 1252
rect 3486 1248 3490 1252
rect 3526 1248 3530 1252
rect 3582 1248 3586 1252
rect 3606 1248 3610 1252
rect 3638 1248 3642 1252
rect 3646 1248 3650 1252
rect 3678 1248 3682 1252
rect 3742 1248 3746 1252
rect 606 1238 610 1242
rect 2838 1238 2842 1242
rect 3198 1238 3202 1242
rect 3622 1238 3626 1242
rect 734 1227 738 1231
rect 838 1227 842 1231
rect 1222 1227 1226 1231
rect 2614 1228 2618 1232
rect 118 1218 122 1222
rect 262 1218 266 1222
rect 446 1218 450 1222
rect 478 1218 482 1222
rect 990 1218 994 1222
rect 1158 1218 1162 1222
rect 1654 1218 1658 1222
rect 1718 1218 1722 1222
rect 1982 1218 1986 1222
rect 2038 1218 2042 1222
rect 2198 1218 2202 1222
rect 2318 1218 2322 1222
rect 2342 1218 2346 1222
rect 2478 1218 2482 1222
rect 2590 1218 2594 1222
rect 2774 1218 2778 1222
rect 2870 1218 2874 1222
rect 2918 1218 2922 1222
rect 2950 1218 2954 1222
rect 2990 1218 2994 1222
rect 3022 1218 3026 1222
rect 3070 1218 3074 1222
rect 3086 1218 3090 1222
rect 3174 1218 3178 1222
rect 3222 1218 3226 1222
rect 3374 1218 3378 1222
rect 3630 1218 3634 1222
rect 346 1203 350 1207
rect 353 1203 357 1207
rect 1362 1203 1366 1207
rect 1369 1203 1373 1207
rect 2386 1203 2390 1207
rect 2393 1203 2397 1207
rect 3410 1203 3414 1207
rect 3417 1203 3421 1207
rect 222 1188 226 1192
rect 246 1188 250 1192
rect 462 1188 466 1192
rect 510 1188 514 1192
rect 598 1188 602 1192
rect 1006 1188 1010 1192
rect 1054 1188 1058 1192
rect 1086 1188 1090 1192
rect 1166 1188 1170 1192
rect 1742 1188 1746 1192
rect 1758 1188 1762 1192
rect 1822 1188 1826 1192
rect 1854 1188 1858 1192
rect 1942 1188 1946 1192
rect 2262 1188 2266 1192
rect 2302 1188 2306 1192
rect 2454 1188 2458 1192
rect 2622 1188 2626 1192
rect 2646 1188 2650 1192
rect 2790 1188 2794 1192
rect 3102 1188 3106 1192
rect 3222 1188 3226 1192
rect 3286 1188 3290 1192
rect 3366 1188 3370 1192
rect 3486 1188 3490 1192
rect 3614 1188 3618 1192
rect 3750 1188 3754 1192
rect 70 1178 74 1182
rect 710 1178 714 1182
rect 206 1168 210 1172
rect 518 1168 522 1172
rect 534 1168 538 1172
rect 1294 1179 1298 1183
rect 1918 1178 1922 1182
rect 2070 1179 2074 1183
rect 3550 1178 3554 1182
rect 846 1168 850 1172
rect 910 1168 914 1172
rect 1550 1168 1554 1172
rect 3494 1168 3498 1172
rect 3534 1168 3538 1172
rect 3606 1168 3610 1172
rect 3726 1168 3730 1172
rect 3758 1168 3762 1172
rect 14 1158 18 1162
rect 70 1148 74 1152
rect 174 1148 178 1152
rect 262 1158 266 1162
rect 326 1158 330 1162
rect 430 1158 434 1162
rect 478 1158 482 1162
rect 502 1158 506 1162
rect 742 1156 746 1160
rect 830 1158 834 1162
rect 878 1158 882 1162
rect 1014 1158 1018 1162
rect 1294 1156 1298 1160
rect 222 1148 226 1152
rect 262 1148 266 1152
rect 278 1148 282 1152
rect 294 1148 298 1152
rect 342 1148 346 1152
rect 422 1148 426 1152
rect 446 1148 450 1152
rect 510 1148 514 1152
rect 534 1148 538 1152
rect 582 1148 586 1152
rect 710 1148 714 1152
rect 806 1148 810 1152
rect 838 1148 842 1152
rect 870 1148 874 1152
rect 894 1148 898 1152
rect 958 1148 962 1152
rect 990 1148 994 1152
rect 1054 1148 1058 1152
rect 1070 1148 1074 1152
rect 1110 1148 1114 1152
rect 1126 1148 1130 1152
rect 1206 1148 1210 1152
rect 1390 1158 1394 1162
rect 1422 1158 1426 1162
rect 1566 1158 1570 1162
rect 1862 1158 1866 1162
rect 1902 1158 1906 1162
rect 1406 1148 1410 1152
rect 1446 1148 1450 1152
rect 1494 1148 1498 1152
rect 1534 1148 1538 1152
rect 1550 1148 1554 1152
rect 1566 1148 1570 1152
rect 1614 1148 1618 1152
rect 1646 1148 1650 1152
rect 1758 1148 1762 1152
rect 1806 1148 1810 1152
rect 2070 1156 2074 1160
rect 2262 1158 2266 1162
rect 2286 1158 2290 1162
rect 2350 1158 2354 1162
rect 2494 1158 2498 1162
rect 2502 1158 2506 1162
rect 2790 1158 2794 1162
rect 2838 1158 2842 1162
rect 1918 1148 1922 1152
rect 2086 1148 2090 1152
rect 2214 1148 2218 1152
rect 2302 1148 2306 1152
rect 2318 1148 2322 1152
rect 2366 1148 2370 1152
rect 2414 1148 2418 1152
rect 2438 1148 2442 1152
rect 2478 1148 2482 1152
rect 2518 1148 2522 1152
rect 2534 1148 2538 1152
rect 2614 1148 2618 1152
rect 2686 1148 2690 1152
rect 2822 1148 2826 1152
rect 2878 1158 2882 1162
rect 2918 1158 2922 1162
rect 2950 1158 2954 1162
rect 3062 1158 3066 1162
rect 3118 1158 3122 1162
rect 3150 1158 3154 1162
rect 3318 1158 3322 1162
rect 3478 1158 3482 1162
rect 3502 1158 3506 1162
rect 3566 1158 3570 1162
rect 3590 1158 3594 1162
rect 3622 1158 3626 1162
rect 3646 1158 3650 1162
rect 3742 1158 3746 1162
rect 3774 1158 3778 1162
rect 2862 1148 2866 1152
rect 2902 1148 2906 1152
rect 2966 1148 2970 1152
rect 2998 1148 3002 1152
rect 3046 1148 3050 1152
rect 3086 1148 3090 1152
rect 3102 1148 3106 1152
rect 3134 1148 3138 1152
rect 3158 1148 3162 1152
rect 3206 1148 3210 1152
rect 3230 1148 3234 1152
rect 3238 1148 3242 1152
rect 3246 1148 3250 1152
rect 3342 1148 3346 1152
rect 3350 1148 3354 1152
rect 3374 1148 3378 1152
rect 3406 1148 3410 1152
rect 3446 1148 3450 1152
rect 3462 1148 3466 1152
rect 3478 1148 3482 1152
rect 3494 1148 3498 1152
rect 3534 1148 3538 1152
rect 3542 1148 3546 1152
rect 3566 1148 3570 1152
rect 3614 1148 3618 1152
rect 3678 1148 3682 1152
rect 3686 1148 3690 1152
rect 3726 1148 3730 1152
rect 3766 1148 3770 1152
rect 70 1138 74 1142
rect 286 1138 290 1142
rect 302 1138 306 1142
rect 334 1138 338 1142
rect 358 1138 362 1142
rect 422 1138 426 1142
rect 438 1138 442 1142
rect 454 1138 458 1142
rect 470 1138 474 1142
rect 494 1138 498 1142
rect 558 1138 562 1142
rect 590 1138 594 1142
rect 710 1138 714 1142
rect 782 1138 786 1142
rect 798 1138 802 1142
rect 902 1138 906 1142
rect 910 1138 914 1142
rect 926 1138 930 1142
rect 998 1138 1002 1142
rect 1038 1138 1042 1142
rect 1046 1138 1050 1142
rect 1078 1138 1082 1142
rect 1102 1138 1106 1142
rect 1262 1138 1266 1142
rect 1334 1138 1338 1142
rect 1350 1138 1354 1142
rect 1414 1138 1418 1142
rect 1438 1138 1442 1142
rect 1494 1138 1498 1142
rect 1518 1138 1522 1142
rect 1558 1138 1562 1142
rect 1606 1138 1610 1142
rect 1638 1138 1642 1142
rect 1686 1138 1690 1142
rect 1798 1138 1802 1142
rect 1814 1138 1818 1142
rect 1862 1138 1866 1142
rect 1878 1138 1882 1142
rect 1926 1138 1930 1142
rect 2038 1138 2042 1142
rect 2214 1138 2218 1142
rect 2310 1138 2314 1142
rect 2326 1138 2330 1142
rect 2374 1138 2378 1142
rect 2382 1138 2386 1142
rect 2398 1138 2402 1142
rect 2462 1138 2466 1142
rect 2470 1138 2474 1142
rect 2510 1138 2514 1142
rect 2526 1138 2530 1142
rect 2542 1138 2546 1142
rect 2574 1138 2578 1142
rect 2742 1138 2746 1142
rect 2814 1138 2818 1142
rect 2846 1138 2850 1142
rect 2870 1138 2874 1142
rect 2894 1138 2898 1142
rect 2942 1138 2946 1142
rect 2982 1138 2986 1142
rect 3006 1138 3010 1142
rect 3014 1138 3018 1142
rect 3038 1138 3042 1142
rect 3054 1138 3058 1142
rect 3094 1138 3098 1142
rect 3126 1138 3130 1142
rect 3254 1138 3258 1142
rect 3286 1138 3290 1142
rect 3302 1138 3306 1142
rect 3334 1138 3338 1142
rect 3454 1138 3458 1142
rect 3542 1138 3546 1142
rect 3574 1138 3578 1142
rect 3630 1138 3634 1142
rect 3646 1138 3650 1142
rect 3710 1138 3714 1142
rect 86 1128 90 1132
rect 238 1128 242 1132
rect 254 1128 258 1132
rect 310 1128 314 1132
rect 318 1128 322 1132
rect 550 1128 554 1132
rect 694 1128 698 1132
rect 1094 1128 1098 1132
rect 1158 1128 1162 1132
rect 1246 1128 1250 1132
rect 1342 1128 1346 1132
rect 1462 1128 1466 1132
rect 1478 1128 1482 1132
rect 1534 1128 1538 1132
rect 1590 1128 1594 1132
rect 1622 1128 1626 1132
rect 1638 1128 1642 1132
rect 1774 1128 1778 1132
rect 1782 1128 1786 1132
rect 2022 1128 2026 1132
rect 2198 1128 2202 1132
rect 2422 1128 2426 1132
rect 2454 1128 2458 1132
rect 2558 1128 2562 1132
rect 2598 1128 2602 1132
rect 2638 1128 2642 1132
rect 2726 1128 2730 1132
rect 2982 1128 2986 1132
rect 3030 1128 3034 1132
rect 3070 1128 3074 1132
rect 3086 1128 3090 1132
rect 3158 1128 3162 1132
rect 3166 1128 3170 1132
rect 3190 1128 3194 1132
rect 3270 1128 3274 1132
rect 3390 1128 3394 1132
rect 3414 1128 3418 1132
rect 3430 1128 3434 1132
rect 3446 1128 3450 1132
rect 3518 1128 3522 1132
rect 190 1118 194 1122
rect 246 1118 250 1122
rect 462 1118 466 1122
rect 486 1118 490 1122
rect 614 1118 618 1122
rect 822 1118 826 1122
rect 942 1118 946 1122
rect 974 1118 978 1122
rect 1006 1118 1010 1122
rect 1030 1118 1034 1122
rect 1126 1118 1130 1122
rect 1382 1118 1386 1122
rect 1430 1118 1434 1122
rect 1670 1118 1674 1122
rect 1766 1118 1770 1122
rect 1790 1118 1794 1122
rect 1822 1118 1826 1122
rect 1942 1118 1946 1122
rect 2118 1118 2122 1122
rect 2334 1118 2338 1122
rect 2494 1118 2498 1122
rect 2582 1118 2586 1122
rect 2886 1118 2890 1122
rect 3022 1118 3026 1122
rect 3646 1118 3650 1122
rect 3702 1118 3706 1122
rect 850 1103 854 1107
rect 857 1103 861 1107
rect 1882 1103 1886 1107
rect 1889 1103 1893 1107
rect 2906 1103 2910 1107
rect 2913 1103 2917 1107
rect 278 1088 282 1092
rect 358 1088 362 1092
rect 742 1088 746 1092
rect 1166 1088 1170 1092
rect 1278 1088 1282 1092
rect 1574 1088 1578 1092
rect 1598 1088 1602 1092
rect 1630 1088 1634 1092
rect 1998 1088 2002 1092
rect 2142 1088 2146 1092
rect 2302 1088 2306 1092
rect 2438 1088 2442 1092
rect 2470 1088 2474 1092
rect 2590 1088 2594 1092
rect 2646 1088 2650 1092
rect 2814 1088 2818 1092
rect 3022 1088 3026 1092
rect 3126 1088 3130 1092
rect 3166 1088 3170 1092
rect 3246 1088 3250 1092
rect 3278 1088 3282 1092
rect 3438 1088 3442 1092
rect 3470 1088 3474 1092
rect 3550 1088 3554 1092
rect 3590 1088 3594 1092
rect 3710 1088 3714 1092
rect 3742 1088 3746 1092
rect 134 1078 138 1082
rect 326 1078 330 1082
rect 438 1078 442 1082
rect 614 1078 618 1082
rect 822 1078 826 1082
rect 998 1078 1002 1082
rect 1470 1078 1474 1082
rect 1510 1078 1514 1082
rect 1526 1078 1530 1082
rect 30 1068 34 1072
rect 118 1068 122 1072
rect 230 1068 234 1072
rect 246 1068 250 1072
rect 454 1068 458 1072
rect 630 1068 634 1072
rect 702 1068 706 1072
rect 838 1068 842 1072
rect 982 1068 986 1072
rect 990 1068 994 1072
rect 1030 1068 1034 1072
rect 1102 1068 1106 1072
rect 1110 1068 1114 1072
rect 1142 1068 1146 1072
rect 1230 1068 1234 1072
rect 1262 1068 1266 1072
rect 1334 1068 1338 1072
rect 1342 1068 1346 1072
rect 1438 1068 1442 1072
rect 1462 1068 1466 1072
rect 1470 1068 1474 1072
rect 1502 1068 1506 1072
rect 1758 1078 1762 1082
rect 1582 1068 1586 1072
rect 1622 1068 1626 1072
rect 1670 1068 1674 1072
rect 1678 1068 1682 1072
rect 1710 1068 1714 1072
rect 1774 1078 1778 1082
rect 1894 1078 1898 1082
rect 2070 1078 2074 1082
rect 2134 1078 2138 1082
rect 2150 1078 2154 1082
rect 2158 1078 2162 1082
rect 2174 1078 2178 1082
rect 2190 1078 2194 1082
rect 2286 1078 2290 1082
rect 1782 1068 1786 1072
rect 1878 1068 1882 1072
rect 2006 1068 2010 1072
rect 2062 1068 2066 1072
rect 2086 1068 2090 1072
rect 2118 1068 2122 1072
rect 2222 1068 2226 1072
rect 2238 1068 2242 1072
rect 2254 1068 2258 1072
rect 2326 1078 2330 1082
rect 2406 1078 2410 1082
rect 2502 1078 2506 1082
rect 2558 1078 2562 1082
rect 2598 1078 2602 1082
rect 2606 1078 2610 1082
rect 2758 1078 2762 1082
rect 2782 1078 2786 1082
rect 2966 1078 2970 1082
rect 3038 1078 3042 1082
rect 3054 1078 3058 1082
rect 3070 1078 3074 1082
rect 3254 1078 3258 1082
rect 3334 1078 3338 1082
rect 3358 1078 3362 1082
rect 3430 1078 3434 1082
rect 3478 1078 3482 1082
rect 3558 1078 3562 1082
rect 2310 1068 2314 1072
rect 2342 1068 2346 1072
rect 2358 1068 2362 1072
rect 2422 1068 2426 1072
rect 2462 1068 2466 1072
rect 2494 1068 2498 1072
rect 2550 1068 2554 1072
rect 2582 1068 2586 1072
rect 2638 1068 2642 1072
rect 2670 1068 2674 1072
rect 2678 1068 2682 1072
rect 2710 1068 2714 1072
rect 2742 1068 2746 1072
rect 2806 1068 2810 1072
rect 2838 1068 2842 1072
rect 2846 1068 2850 1072
rect 2862 1068 2866 1072
rect 2942 1068 2946 1072
rect 3118 1068 3122 1072
rect 3142 1068 3146 1072
rect 3238 1068 3242 1072
rect 3262 1068 3266 1072
rect 3462 1068 3466 1072
rect 3486 1068 3490 1072
rect 3510 1068 3514 1072
rect 3566 1068 3570 1072
rect 3598 1068 3602 1072
rect 3622 1068 3626 1072
rect 3686 1068 3690 1072
rect 3718 1068 3722 1072
rect 22 1058 26 1062
rect 46 1058 50 1062
rect 174 1058 178 1062
rect 262 1058 266 1062
rect 302 1058 306 1062
rect 326 1058 330 1062
rect 398 1058 402 1062
rect 574 1058 578 1062
rect 710 1058 714 1062
rect 726 1058 730 1062
rect 782 1058 786 1062
rect 942 1058 946 1062
rect 958 1058 962 1062
rect 974 1058 978 1062
rect 1014 1058 1018 1062
rect 1022 1058 1026 1062
rect 1118 1058 1122 1062
rect 1134 1058 1138 1062
rect 1150 1058 1154 1062
rect 1190 1058 1194 1062
rect 1214 1058 1218 1062
rect 1222 1058 1226 1062
rect 1238 1058 1242 1062
rect 1254 1058 1258 1062
rect 1374 1058 1378 1062
rect 1390 1058 1394 1062
rect 1398 1058 1402 1062
rect 1494 1058 1498 1062
rect 1510 1058 1514 1062
rect 1534 1058 1538 1062
rect 1590 1058 1594 1062
rect 1638 1058 1642 1062
rect 1662 1058 1666 1062
rect 1686 1058 1690 1062
rect 1718 1058 1722 1062
rect 1742 1058 1746 1062
rect 1798 1058 1802 1062
rect 1830 1058 1834 1062
rect 2014 1058 2018 1062
rect 2054 1058 2058 1062
rect 2094 1058 2098 1062
rect 2174 1058 2178 1062
rect 2198 1058 2202 1062
rect 2230 1058 2234 1062
rect 2246 1058 2250 1062
rect 2262 1058 2266 1062
rect 2270 1058 2274 1062
rect 2350 1058 2354 1062
rect 2358 1058 2362 1062
rect 2430 1058 2434 1062
rect 2454 1058 2458 1062
rect 2486 1058 2490 1062
rect 2518 1058 2522 1062
rect 2526 1058 2530 1062
rect 2542 1058 2546 1062
rect 2574 1058 2578 1062
rect 2614 1058 2618 1062
rect 2630 1058 2634 1062
rect 2662 1058 2666 1062
rect 2686 1058 2690 1062
rect 2718 1058 2722 1062
rect 2734 1058 2738 1062
rect 2766 1058 2770 1062
rect 2774 1058 2778 1062
rect 2790 1058 2794 1062
rect 2806 1058 2810 1062
rect 2830 1058 2834 1062
rect 2918 1058 2922 1062
rect 2934 1058 2938 1062
rect 2950 1058 2954 1062
rect 2974 1058 2978 1062
rect 2998 1058 3002 1062
rect 3054 1058 3058 1062
rect 3094 1058 3098 1062
rect 3110 1058 3114 1062
rect 3142 1058 3146 1062
rect 3150 1058 3154 1062
rect 3182 1058 3186 1062
rect 3214 1058 3218 1062
rect 3222 1058 3226 1062
rect 3230 1058 3234 1062
rect 3286 1058 3290 1062
rect 3294 1058 3298 1062
rect 3318 1058 3322 1062
rect 3358 1058 3362 1062
rect 3382 1058 3386 1062
rect 3390 1058 3394 1062
rect 3446 1058 3450 1062
rect 3454 1058 3458 1062
rect 3502 1058 3506 1062
rect 3534 1058 3538 1062
rect 3574 1058 3578 1062
rect 3622 1058 3626 1062
rect 3630 1058 3634 1062
rect 3678 1058 3682 1062
rect 3694 1058 3698 1062
rect 3726 1058 3730 1062
rect 3774 1058 3778 1062
rect 70 1048 74 1052
rect 254 1048 258 1052
rect 326 1048 330 1052
rect 502 1048 506 1052
rect 678 1048 682 1052
rect 870 1050 874 1054
rect 950 1048 954 1052
rect 958 1048 962 1052
rect 1006 1048 1010 1052
rect 1358 1048 1362 1052
rect 1382 1048 1386 1052
rect 1414 1048 1418 1052
rect 1478 1048 1482 1052
rect 1598 1048 1602 1052
rect 1638 1048 1642 1052
rect 1646 1048 1650 1052
rect 1702 1048 1706 1052
rect 1718 1048 1722 1052
rect 1734 1048 1738 1052
rect 1846 1050 1850 1054
rect 2014 1048 2018 1052
rect 2030 1048 2034 1052
rect 2038 1048 2042 1052
rect 2070 1048 2074 1052
rect 2102 1048 2106 1052
rect 2366 1048 2370 1052
rect 2438 1048 2442 1052
rect 2470 1048 2474 1052
rect 2566 1048 2570 1052
rect 2606 1048 2610 1052
rect 2646 1048 2650 1052
rect 2702 1048 2706 1052
rect 2718 1048 2722 1052
rect 2814 1048 2818 1052
rect 2862 1048 2866 1052
rect 2918 1048 2922 1052
rect 3070 1048 3074 1052
rect 3102 1048 3106 1052
rect 3278 1048 3282 1052
rect 3406 1048 3410 1052
rect 3502 1048 3506 1052
rect 3526 1048 3530 1052
rect 3590 1048 3594 1052
rect 3614 1048 3618 1052
rect 3646 1048 3650 1052
rect 3662 1048 3666 1052
rect 6 1038 10 1042
rect 294 1038 298 1042
rect 310 1038 314 1042
rect 934 1038 938 1042
rect 3094 1038 3098 1042
rect 3350 1038 3354 1042
rect 174 1027 178 1031
rect 398 1027 402 1031
rect 574 1027 578 1031
rect 870 1027 874 1031
rect 2126 1028 2130 1032
rect 2934 1028 2938 1032
rect 3630 1028 3634 1032
rect 214 1018 218 1022
rect 238 1018 242 1022
rect 302 1018 306 1022
rect 534 1018 538 1022
rect 926 1018 930 1022
rect 998 1018 1002 1022
rect 1046 1018 1050 1022
rect 1134 1018 1138 1022
rect 1166 1018 1170 1022
rect 1198 1018 1202 1022
rect 1254 1018 1258 1022
rect 1550 1018 1554 1022
rect 1686 1018 1690 1022
rect 1846 1018 1850 1022
rect 1974 1018 1978 1022
rect 2054 1018 2058 1022
rect 2174 1018 2178 1022
rect 2510 1018 2514 1022
rect 2686 1018 2690 1022
rect 2750 1018 2754 1022
rect 2950 1018 2954 1022
rect 2990 1018 2994 1022
rect 3046 1018 3050 1022
rect 3206 1018 3210 1022
rect 3310 1018 3314 1022
rect 3390 1018 3394 1022
rect 3758 1018 3762 1022
rect 346 1003 350 1007
rect 353 1003 357 1007
rect 1362 1003 1366 1007
rect 1369 1003 1373 1007
rect 2386 1003 2390 1007
rect 2393 1003 2397 1007
rect 3410 1003 3414 1007
rect 3417 1003 3421 1007
rect 14 988 18 992
rect 374 988 378 992
rect 422 988 426 992
rect 454 988 458 992
rect 574 988 578 992
rect 718 988 722 992
rect 758 988 762 992
rect 902 988 906 992
rect 1126 988 1130 992
rect 1238 988 1242 992
rect 1382 988 1386 992
rect 1574 988 1578 992
rect 1790 988 1794 992
rect 2150 988 2154 992
rect 2934 988 2938 992
rect 3550 988 3554 992
rect 3614 988 3618 992
rect 3670 988 3674 992
rect 102 978 106 982
rect 238 978 242 982
rect 998 979 1002 983
rect 1446 978 1450 982
rect 1774 978 1778 982
rect 2022 979 2026 983
rect 2190 978 2194 982
rect 3046 978 3050 982
rect 446 968 450 972
rect 494 968 498 972
rect 2294 968 2298 972
rect 2670 968 2674 972
rect 3038 968 3042 972
rect 3334 968 3338 972
rect 3382 968 3386 972
rect 3486 968 3490 972
rect 3494 968 3498 972
rect 3542 968 3546 972
rect 3574 968 3578 972
rect 3582 968 3586 972
rect 3606 968 3610 972
rect 3662 968 3666 972
rect 46 958 50 962
rect 70 956 74 960
rect 262 958 266 962
rect 286 958 290 962
rect 326 958 330 962
rect 30 948 34 952
rect 102 948 106 952
rect 310 948 314 952
rect 342 948 346 952
rect 390 948 394 952
rect 462 958 466 962
rect 542 958 546 962
rect 718 958 722 962
rect 758 958 762 962
rect 926 958 930 962
rect 998 956 1002 960
rect 1382 958 1386 962
rect 1590 958 1594 962
rect 1630 958 1634 962
rect 1678 958 1682 962
rect 454 948 458 952
rect 470 948 474 952
rect 702 948 706 952
rect 758 948 762 952
rect 918 948 922 952
rect 950 948 954 952
rect 1086 948 1090 952
rect 1142 948 1146 952
rect 1158 948 1162 952
rect 1174 948 1178 952
rect 1206 948 1210 952
rect 1278 948 1282 952
rect 1374 948 1378 952
rect 1438 948 1442 952
rect 1558 948 1562 952
rect 1574 948 1578 952
rect 1598 948 1602 952
rect 1654 948 1658 952
rect 1710 958 1714 962
rect 1926 958 1930 962
rect 2022 956 2026 960
rect 2222 958 2226 962
rect 2246 958 2250 962
rect 2278 958 2282 962
rect 2302 958 2306 962
rect 2334 958 2338 962
rect 2366 958 2370 962
rect 2478 958 2482 962
rect 2558 958 2562 962
rect 2566 958 2570 962
rect 2638 958 2642 962
rect 2654 958 2658 962
rect 2726 958 2730 962
rect 2798 958 2802 962
rect 2814 958 2818 962
rect 2830 958 2834 962
rect 2902 958 2906 962
rect 2950 958 2954 962
rect 2958 958 2962 962
rect 3014 958 3018 962
rect 3078 958 3082 962
rect 3142 958 3146 962
rect 3150 958 3154 962
rect 3206 958 3210 962
rect 3262 958 3266 962
rect 3366 958 3370 962
rect 3398 958 3402 962
rect 3470 958 3474 962
rect 3502 958 3506 962
rect 3558 958 3562 962
rect 3590 958 3594 962
rect 3622 958 3626 962
rect 3646 958 3650 962
rect 3678 958 3682 962
rect 3710 958 3714 962
rect 3774 958 3778 962
rect 1726 948 1730 952
rect 1742 948 1746 952
rect 1822 948 1826 952
rect 1854 948 1858 952
rect 1878 948 1882 952
rect 1910 948 1914 952
rect 1958 948 1962 952
rect 2110 948 2114 952
rect 2166 948 2170 952
rect 2198 948 2202 952
rect 2262 948 2266 952
rect 2278 948 2282 952
rect 2310 948 2314 952
rect 2382 948 2386 952
rect 2414 948 2418 952
rect 2470 948 2474 952
rect 2494 948 2498 952
rect 2526 948 2530 952
rect 2542 948 2546 952
rect 2582 948 2586 952
rect 2590 948 2594 952
rect 2630 948 2634 952
rect 2718 948 2722 952
rect 2742 948 2746 952
rect 2774 948 2778 952
rect 2806 948 2810 952
rect 102 938 106 942
rect 230 938 234 942
rect 262 938 266 942
rect 302 938 306 942
rect 430 938 434 942
rect 470 938 474 942
rect 494 938 498 942
rect 526 938 530 942
rect 566 938 570 942
rect 670 938 674 942
rect 806 938 810 942
rect 958 938 962 942
rect 1030 938 1034 942
rect 1150 938 1154 942
rect 1334 938 1338 942
rect 1526 938 1530 942
rect 1550 938 1554 942
rect 1566 938 1570 942
rect 1606 938 1610 942
rect 1622 938 1626 942
rect 1654 938 1658 942
rect 1662 938 1666 942
rect 1686 938 1690 942
rect 1734 938 1738 942
rect 1766 938 1770 942
rect 1782 938 1786 942
rect 1830 938 1834 942
rect 1846 938 1850 942
rect 1894 938 1898 942
rect 2054 938 2058 942
rect 2174 938 2178 942
rect 2190 938 2194 942
rect 2206 938 2210 942
rect 2222 938 2226 942
rect 2230 938 2234 942
rect 2254 938 2258 942
rect 2286 938 2290 942
rect 2326 938 2330 942
rect 2358 938 2362 942
rect 2390 938 2394 942
rect 2446 938 2450 942
rect 2462 938 2466 942
rect 2502 938 2506 942
rect 2534 938 2538 942
rect 2574 938 2578 942
rect 2590 938 2594 942
rect 2606 938 2610 942
rect 2670 938 2674 942
rect 2686 938 2690 942
rect 2758 938 2762 942
rect 2782 938 2786 942
rect 2798 938 2802 942
rect 2838 948 2842 952
rect 2870 948 2874 952
rect 2886 948 2890 952
rect 2918 948 2922 952
rect 2934 948 2938 952
rect 2974 948 2978 952
rect 2998 948 3002 952
rect 3030 948 3034 952
rect 3062 948 3066 952
rect 3070 948 3074 952
rect 3086 948 3090 952
rect 3126 948 3130 952
rect 3230 948 3234 952
rect 3246 948 3250 952
rect 3286 948 3290 952
rect 3310 948 3314 952
rect 3334 948 3338 952
rect 3342 948 3346 952
rect 3366 948 3370 952
rect 3390 948 3394 952
rect 3406 948 3410 952
rect 3494 948 3498 952
rect 3526 948 3530 952
rect 3550 948 3554 952
rect 3582 948 3586 952
rect 3614 948 3618 952
rect 3670 948 3674 952
rect 3686 948 3690 952
rect 3726 948 3730 952
rect 3766 948 3770 952
rect 2846 938 2850 942
rect 2862 938 2866 942
rect 2878 938 2882 942
rect 2926 938 2930 942
rect 2982 938 2986 942
rect 2990 938 2994 942
rect 3054 938 3058 942
rect 3094 938 3098 942
rect 3118 938 3122 942
rect 3134 938 3138 942
rect 3166 938 3170 942
rect 3182 938 3186 942
rect 3190 938 3194 942
rect 3238 938 3242 942
rect 3286 938 3290 942
rect 3294 938 3298 942
rect 3342 938 3346 942
rect 3382 938 3386 942
rect 3446 938 3450 942
rect 3630 938 3634 942
rect 3686 938 3690 942
rect 3750 938 3754 942
rect 118 928 122 932
rect 214 928 218 932
rect 406 928 410 932
rect 534 928 538 932
rect 566 928 570 932
rect 654 928 658 932
rect 822 928 826 932
rect 1046 928 1050 932
rect 1182 928 1186 932
rect 1222 928 1226 932
rect 1318 928 1322 932
rect 1422 928 1426 932
rect 1454 928 1458 932
rect 1534 928 1538 932
rect 1622 928 1626 932
rect 1798 928 1802 932
rect 1806 928 1810 932
rect 1814 928 1818 932
rect 1838 928 1842 932
rect 1862 928 1866 932
rect 1950 928 1954 932
rect 1974 928 1978 932
rect 2070 928 2074 932
rect 2446 928 2450 932
rect 2478 928 2482 932
rect 2510 928 2514 932
rect 2622 928 2626 932
rect 2646 928 2650 932
rect 2846 928 2850 932
rect 3110 928 3114 932
rect 3174 928 3178 932
rect 3214 928 3218 932
rect 3270 928 3274 932
rect 3294 928 3298 932
rect 3318 928 3322 932
rect 3422 928 3426 932
rect 3510 928 3514 932
rect 14 918 18 922
rect 198 918 202 922
rect 270 918 274 922
rect 286 918 290 922
rect 550 918 554 922
rect 1430 918 1434 922
rect 1470 918 1474 922
rect 1542 918 1546 922
rect 1614 918 1618 922
rect 1670 918 1674 922
rect 1702 918 1706 922
rect 1870 918 1874 922
rect 1926 918 1930 922
rect 1942 918 1946 922
rect 2246 918 2250 922
rect 2430 918 2434 922
rect 2518 918 2522 922
rect 2558 918 2562 922
rect 2614 918 2618 922
rect 2662 918 2666 922
rect 2702 918 2706 922
rect 2726 918 2730 922
rect 2766 918 2770 922
rect 2830 918 2834 922
rect 2958 918 2962 922
rect 3102 918 3106 922
rect 3150 918 3154 922
rect 3206 918 3210 922
rect 3262 918 3266 922
rect 3470 918 3474 922
rect 3518 918 3522 922
rect 3638 918 3642 922
rect 850 903 854 907
rect 857 903 861 907
rect 1882 903 1886 907
rect 1889 903 1893 907
rect 2906 903 2910 907
rect 2913 903 2917 907
rect 222 888 226 892
rect 238 888 242 892
rect 438 888 442 892
rect 534 888 538 892
rect 926 888 930 892
rect 1174 888 1178 892
rect 1294 888 1298 892
rect 1606 888 1610 892
rect 1862 888 1866 892
rect 1918 888 1922 892
rect 1958 888 1962 892
rect 2374 888 2378 892
rect 2398 888 2402 892
rect 2446 888 2450 892
rect 2550 888 2554 892
rect 3374 888 3378 892
rect 3590 888 3594 892
rect 3718 888 3722 892
rect 86 878 90 882
rect 182 878 186 882
rect 310 878 314 882
rect 334 878 338 882
rect 366 878 370 882
rect 414 878 418 882
rect 462 878 466 882
rect 542 878 546 882
rect 590 878 594 882
rect 742 878 746 882
rect 1006 878 1010 882
rect 1142 878 1146 882
rect 1198 878 1202 882
rect 1254 878 1258 882
rect 1286 878 1290 882
rect 1310 878 1314 882
rect 1414 878 1418 882
rect 1638 878 1642 882
rect 1710 878 1714 882
rect 1766 878 1770 882
rect 1902 878 1906 882
rect 2038 878 2042 882
rect 2214 878 2218 882
rect 2334 878 2338 882
rect 2438 878 2442 882
rect 2470 878 2474 882
rect 2486 878 2490 882
rect 2510 878 2514 882
rect 2518 878 2522 882
rect 2542 878 2546 882
rect 2566 878 2570 882
rect 2678 878 2682 882
rect 2878 878 2882 882
rect 2926 878 2930 882
rect 3030 878 3034 882
rect 3038 878 3042 882
rect 3206 878 3210 882
rect 3270 878 3274 882
rect 3278 878 3282 882
rect 3302 878 3306 882
rect 3326 878 3330 882
rect 3382 878 3386 882
rect 3406 878 3410 882
rect 3526 878 3530 882
rect 70 868 74 872
rect 198 868 202 872
rect 294 868 298 872
rect 398 868 402 872
rect 430 868 434 872
rect 446 868 450 872
rect 478 868 482 872
rect 510 868 514 872
rect 550 868 554 872
rect 646 868 650 872
rect 758 868 762 872
rect 846 868 850 872
rect 1022 868 1026 872
rect 1158 868 1162 872
rect 1190 868 1194 872
rect 1214 868 1218 872
rect 1230 868 1234 872
rect 1278 868 1282 872
rect 1430 868 1434 872
rect 1502 868 1506 872
rect 1558 868 1562 872
rect 1582 868 1586 872
rect 1598 868 1602 872
rect 1742 868 1746 872
rect 1774 868 1778 872
rect 1846 868 1850 872
rect 1862 868 1866 872
rect 1902 868 1906 872
rect 1950 868 1954 872
rect 2054 868 2058 872
rect 2230 868 2234 872
rect 2302 868 2306 872
rect 2358 868 2362 872
rect 2366 868 2370 872
rect 2430 868 2434 872
rect 2454 868 2458 872
rect 2590 868 2594 872
rect 2606 868 2610 872
rect 2622 868 2626 872
rect 2638 868 2642 872
rect 2662 868 2666 872
rect 2686 868 2690 872
rect 2742 868 2746 872
rect 2750 868 2754 872
rect 2766 868 2770 872
rect 2782 868 2786 872
rect 2798 868 2802 872
rect 2814 868 2818 872
rect 2846 868 2850 872
rect 2894 868 2898 872
rect 2942 868 2946 872
rect 2958 868 2962 872
rect 2990 868 2994 872
rect 3014 868 3018 872
rect 3022 868 3026 872
rect 3046 868 3050 872
rect 3094 868 3098 872
rect 3126 868 3130 872
rect 3134 868 3138 872
rect 3166 868 3170 872
rect 3206 868 3210 872
rect 3246 868 3250 872
rect 3254 868 3258 872
rect 3270 868 3274 872
rect 3318 868 3322 872
rect 3350 868 3354 872
rect 3398 868 3402 872
rect 3462 868 3466 872
rect 3478 868 3482 872
rect 3502 868 3506 872
rect 3518 868 3522 872
rect 3558 868 3562 872
rect 3630 868 3634 872
rect 3694 868 3698 872
rect 3726 868 3730 872
rect 126 858 130 862
rect 318 858 322 862
rect 382 858 386 862
rect 390 858 394 862
rect 406 858 410 862
rect 422 858 426 862
rect 454 858 458 862
rect 486 858 490 862
rect 502 858 506 862
rect 558 858 562 862
rect 702 858 706 862
rect 910 858 914 862
rect 1070 858 1074 862
rect 1102 858 1106 862
rect 1126 858 1130 862
rect 1134 858 1138 862
rect 1166 858 1170 862
rect 1206 858 1210 862
rect 1222 858 1226 862
rect 1278 858 1282 862
rect 1302 858 1306 862
rect 1374 858 1378 862
rect 1478 858 1482 862
rect 1510 858 1514 862
rect 1534 858 1538 862
rect 1550 858 1554 862
rect 1590 858 1594 862
rect 1622 858 1626 862
rect 1662 858 1666 862
rect 1678 858 1682 862
rect 1710 858 1714 862
rect 1734 858 1738 862
rect 1750 858 1754 862
rect 1782 858 1786 862
rect 1830 858 1834 862
rect 1838 858 1842 862
rect 1870 858 1874 862
rect 1910 858 1914 862
rect 1942 858 1946 862
rect 1998 858 2002 862
rect 2110 858 2114 862
rect 2174 858 2178 862
rect 2286 858 2290 862
rect 2310 858 2314 862
rect 2350 858 2354 862
rect 2422 858 2426 862
rect 2462 858 2466 862
rect 2494 858 2498 862
rect 2534 858 2538 862
rect 2558 858 2562 862
rect 2582 858 2586 862
rect 2614 858 2618 862
rect 2630 858 2634 862
rect 2654 858 2658 862
rect 2670 858 2674 862
rect 2686 858 2690 862
rect 2734 858 2738 862
rect 2774 858 2778 862
rect 2806 858 2810 862
rect 2822 858 2826 862
rect 2854 858 2858 862
rect 2902 858 2906 862
rect 2950 858 2954 862
rect 2974 858 2978 862
rect 2982 858 2986 862
rect 3086 858 3090 862
rect 3118 858 3122 862
rect 3142 858 3146 862
rect 3174 858 3178 862
rect 3230 858 3234 862
rect 3238 858 3242 862
rect 3294 858 3298 862
rect 3318 858 3322 862
rect 3342 858 3346 862
rect 3358 858 3362 862
rect 3398 858 3402 862
rect 3454 858 3458 862
rect 3470 858 3474 862
rect 3510 858 3514 862
rect 3558 858 3562 862
rect 3574 858 3578 862
rect 3630 858 3634 862
rect 3638 858 3642 862
rect 3662 858 3666 862
rect 3686 858 3690 862
rect 3702 858 3706 862
rect 3750 858 3754 862
rect 14 848 18 852
rect 222 848 226 852
rect 574 848 578 852
rect 790 850 794 854
rect 1054 850 1058 854
rect 1174 848 1178 852
rect 1462 850 1466 854
rect 1510 848 1514 852
rect 1526 848 1530 852
rect 1534 848 1538 852
rect 1566 848 1570 852
rect 1646 848 1650 852
rect 1718 848 1722 852
rect 1782 848 1786 852
rect 1798 848 1802 852
rect 1886 848 1890 852
rect 2102 848 2106 852
rect 2262 850 2266 854
rect 2326 848 2330 852
rect 2382 848 2386 852
rect 2390 848 2394 852
rect 2646 848 2650 852
rect 2710 848 2714 852
rect 2766 848 2770 852
rect 2838 848 2842 852
rect 2934 848 2938 852
rect 2966 848 2970 852
rect 2998 848 3002 852
rect 3070 848 3074 852
rect 3102 848 3106 852
rect 3118 848 3122 852
rect 3158 848 3162 852
rect 3190 848 3194 852
rect 3214 848 3218 852
rect 3374 848 3378 852
rect 3486 848 3490 852
rect 3494 848 3498 852
rect 3590 848 3594 852
rect 3654 848 3658 852
rect 382 838 386 842
rect 2798 838 2802 842
rect 3174 838 3178 842
rect 3342 838 3346 842
rect 3454 838 3458 842
rect 3558 838 3562 842
rect 126 827 130 831
rect 790 827 794 831
rect 1054 827 1058 831
rect 1462 827 1466 831
rect 1662 828 1666 832
rect 2262 827 2266 831
rect 3086 828 3090 832
rect 3606 828 3610 832
rect 166 818 170 822
rect 302 818 306 822
rect 470 818 474 822
rect 558 818 562 822
rect 662 818 666 822
rect 1118 818 1122 822
rect 1142 818 1146 822
rect 1238 818 1242 822
rect 1814 818 1818 822
rect 2102 818 2106 822
rect 2134 818 2138 822
rect 2478 818 2482 822
rect 2526 818 2530 822
rect 2550 818 2554 822
rect 2694 818 2698 822
rect 2734 818 2738 822
rect 2822 818 2826 822
rect 2854 818 2858 822
rect 3006 818 3010 822
rect 3062 818 3066 822
rect 3142 818 3146 822
rect 3230 818 3234 822
rect 3294 818 3298 822
rect 3670 818 3674 822
rect 346 803 350 807
rect 353 803 357 807
rect 1362 803 1366 807
rect 1369 803 1373 807
rect 2386 803 2390 807
rect 2393 803 2397 807
rect 3410 803 3414 807
rect 3417 803 3421 807
rect 278 788 282 792
rect 390 788 394 792
rect 494 788 498 792
rect 790 788 794 792
rect 902 788 906 792
rect 1126 788 1130 792
rect 1326 788 1330 792
rect 1470 788 1474 792
rect 1782 788 1786 792
rect 1846 788 1850 792
rect 2342 788 2346 792
rect 2366 788 2370 792
rect 2494 788 2498 792
rect 2518 788 2522 792
rect 2662 788 2666 792
rect 3134 788 3138 792
rect 3430 788 3434 792
rect 3518 788 3522 792
rect 3542 788 3546 792
rect 3582 788 3586 792
rect 3614 788 3618 792
rect 190 778 194 782
rect 638 778 642 782
rect 318 768 322 772
rect 366 768 370 772
rect 998 779 1002 783
rect 1686 778 1690 782
rect 2022 779 2026 783
rect 830 768 834 772
rect 1894 768 1898 772
rect 2862 768 2866 772
rect 3094 768 3098 772
rect 3190 768 3194 772
rect 3550 768 3554 772
rect 3622 768 3626 772
rect 3670 768 3674 772
rect 3710 768 3714 772
rect 3726 768 3730 772
rect 3758 768 3762 772
rect 54 758 58 762
rect 174 758 178 762
rect 294 758 298 762
rect 302 758 306 762
rect 462 758 466 762
rect 486 758 490 762
rect 670 756 674 760
rect 814 758 818 762
rect 998 756 1002 760
rect 1142 758 1146 762
rect 1206 758 1210 762
rect 1222 758 1226 762
rect 1470 758 1474 762
rect 1542 758 1546 762
rect 1574 758 1578 762
rect 1630 758 1634 762
rect 1702 758 1706 762
rect 30 748 34 752
rect 70 748 74 752
rect 166 748 170 752
rect 190 748 194 752
rect 206 748 210 752
rect 262 748 266 752
rect 278 748 282 752
rect 358 748 362 752
rect 398 748 402 752
rect 406 748 410 752
rect 446 748 450 752
rect 502 748 506 752
rect 510 748 514 752
rect 638 748 642 752
rect 790 748 794 752
rect 822 748 826 752
rect 862 748 866 752
rect 1086 748 1090 752
rect 1166 748 1170 752
rect 1182 748 1186 752
rect 2022 756 2026 760
rect 2078 758 2082 762
rect 1254 748 1258 752
rect 1294 748 1298 752
rect 1478 748 1482 752
rect 1510 748 1514 752
rect 1518 748 1522 752
rect 1558 748 1562 752
rect 1566 748 1570 752
rect 1614 748 1618 752
rect 1630 748 1634 752
rect 1670 748 1674 752
rect 1686 748 1690 752
rect 1726 748 1730 752
rect 1734 748 1738 752
rect 1766 748 1770 752
rect 1798 748 1802 752
rect 1806 748 1810 752
rect 1830 748 1834 752
rect 1862 748 1866 752
rect 1934 748 1938 752
rect 2214 758 2218 762
rect 2358 758 2362 762
rect 2430 758 2434 762
rect 2518 758 2522 762
rect 2910 758 2914 762
rect 2974 758 2978 762
rect 3078 758 3082 762
rect 3166 758 3170 762
rect 3254 758 3258 762
rect 3374 758 3378 762
rect 3446 758 3450 762
rect 3462 758 3466 762
rect 3502 758 3506 762
rect 3534 758 3538 762
rect 3566 758 3570 762
rect 3598 758 3602 762
rect 3606 758 3610 762
rect 3654 758 3658 762
rect 3686 758 3690 762
rect 3742 758 3746 762
rect 3774 758 3778 762
rect 2102 748 2106 752
rect 2134 748 2138 752
rect 2174 748 2178 752
rect 2206 748 2210 752
rect 2238 748 2242 752
rect 2262 748 2266 752
rect 2318 748 2322 752
rect 2342 748 2346 752
rect 2422 748 2426 752
rect 2446 748 2450 752
rect 2454 748 2458 752
rect 2486 748 2490 752
rect 2518 748 2522 752
rect 2702 748 2706 752
rect 2734 748 2738 752
rect 2750 748 2754 752
rect 2766 748 2770 752
rect 2798 748 2802 752
rect 2822 748 2826 752
rect 2830 748 2834 752
rect 2886 748 2890 752
rect 2926 748 2930 752
rect 2958 748 2962 752
rect 2974 748 2978 752
rect 3022 748 3026 752
rect 3030 748 3034 752
rect 3110 748 3114 752
rect 3142 748 3146 752
rect 3190 748 3194 752
rect 78 738 82 742
rect 94 738 98 742
rect 134 738 138 742
rect 142 738 146 742
rect 158 738 162 742
rect 198 738 202 742
rect 214 738 218 742
rect 238 738 242 742
rect 254 738 258 742
rect 270 738 274 742
rect 454 738 458 742
rect 478 738 482 742
rect 638 738 642 742
rect 774 738 778 742
rect 782 738 786 742
rect 894 738 898 742
rect 958 738 962 742
rect 1030 738 1034 742
rect 1158 738 1162 742
rect 1174 738 1178 742
rect 1190 738 1194 742
rect 1222 738 1226 742
rect 1422 738 1426 742
rect 1510 738 1514 742
rect 1550 738 1554 742
rect 1606 738 1610 742
rect 1742 738 1746 742
rect 1774 738 1778 742
rect 1990 738 1994 742
rect 2062 738 2066 742
rect 2078 738 2082 742
rect 2110 738 2114 742
rect 2142 738 2146 742
rect 2150 738 2154 742
rect 2166 738 2170 742
rect 2230 738 2234 742
rect 2294 738 2298 742
rect 2326 738 2330 742
rect 2334 738 2338 742
rect 2414 738 2418 742
rect 2438 738 2442 742
rect 2454 738 2458 742
rect 2486 738 2490 742
rect 2566 738 2570 742
rect 2694 738 2698 742
rect 2726 738 2730 742
rect 2742 738 2746 742
rect 2798 738 2802 742
rect 2838 738 2842 742
rect 2878 738 2882 742
rect 2934 738 2938 742
rect 2966 738 2970 742
rect 3014 738 3018 742
rect 3102 738 3106 742
rect 3118 738 3122 742
rect 3134 738 3138 742
rect 3238 748 3242 752
rect 3262 748 3266 752
rect 3286 748 3290 752
rect 3326 748 3330 752
rect 3342 748 3346 752
rect 3358 748 3362 752
rect 3382 748 3386 752
rect 3398 748 3402 752
rect 3478 748 3482 752
rect 3486 748 3490 752
rect 3518 748 3522 752
rect 3558 748 3562 752
rect 3582 748 3586 752
rect 3614 748 3618 752
rect 3678 748 3682 752
rect 3710 748 3714 752
rect 3718 748 3722 752
rect 3766 748 3770 752
rect 3206 738 3210 742
rect 3230 738 3234 742
rect 3246 738 3250 742
rect 3302 738 3306 742
rect 3350 738 3354 742
rect 3422 738 3426 742
rect 3478 738 3482 742
rect 3510 738 3514 742
rect 3574 738 3578 742
rect 3638 738 3642 742
rect 3654 738 3658 742
rect 3678 738 3682 742
rect 3718 738 3722 742
rect 134 728 138 732
rect 142 728 146 732
rect 230 728 234 732
rect 238 728 242 732
rect 334 728 338 732
rect 382 728 386 732
rect 422 728 426 732
rect 462 728 466 732
rect 526 728 530 732
rect 622 728 626 732
rect 1046 728 1050 732
rect 1230 728 1234 732
rect 1270 728 1274 732
rect 1278 728 1282 732
rect 1406 728 1410 732
rect 1494 728 1498 732
rect 1598 728 1602 732
rect 1638 728 1642 732
rect 1710 728 1714 732
rect 1974 728 1978 732
rect 2150 728 2154 732
rect 2190 728 2194 732
rect 2374 728 2378 732
rect 2398 728 2402 732
rect 2478 728 2482 732
rect 2582 728 2586 732
rect 2678 728 2682 732
rect 2710 728 2714 732
rect 2718 728 2722 732
rect 2774 728 2778 732
rect 2806 728 2810 732
rect 2854 728 2858 732
rect 2862 728 2866 732
rect 2942 728 2946 732
rect 2958 728 2962 732
rect 2998 728 3002 732
rect 3046 728 3050 732
rect 3054 728 3058 732
rect 3086 728 3090 732
rect 3134 728 3138 732
rect 3174 728 3178 732
rect 3222 728 3226 732
rect 3278 728 3282 732
rect 3302 728 3306 732
rect 3310 728 3314 732
rect 3326 728 3330 732
rect 3382 728 3386 732
rect 3454 728 3458 732
rect 3502 728 3506 732
rect 3694 728 3698 732
rect 14 718 18 722
rect 86 718 90 722
rect 222 718 226 722
rect 414 718 418 722
rect 430 718 434 722
rect 718 718 722 722
rect 878 718 882 722
rect 1142 718 1146 722
rect 1502 718 1506 722
rect 1542 718 1546 722
rect 1718 718 1722 722
rect 1750 718 1754 722
rect 1846 718 1850 722
rect 2118 718 2122 722
rect 2214 718 2218 722
rect 2254 718 2258 722
rect 2302 718 2306 722
rect 2366 718 2370 722
rect 2406 718 2410 722
rect 2662 718 2666 722
rect 2686 718 2690 722
rect 2814 718 2818 722
rect 2846 718 2850 722
rect 2894 718 2898 722
rect 3038 718 3042 722
rect 3062 718 3066 722
rect 3166 718 3170 722
rect 3214 718 3218 722
rect 3270 718 3274 722
rect 3318 718 3322 722
rect 3750 718 3754 722
rect 850 703 854 707
rect 857 703 861 707
rect 1882 703 1886 707
rect 1889 703 1893 707
rect 2906 703 2910 707
rect 2913 703 2917 707
rect 270 688 274 692
rect 294 688 298 692
rect 390 688 394 692
rect 550 688 554 692
rect 606 688 610 692
rect 830 688 834 692
rect 886 688 890 692
rect 1502 688 1506 692
rect 1958 688 1962 692
rect 2054 688 2058 692
rect 2454 688 2458 692
rect 2486 688 2490 692
rect 2542 688 2546 692
rect 2798 688 2802 692
rect 2838 688 2842 692
rect 2870 688 2874 692
rect 2902 688 2906 692
rect 2982 688 2986 692
rect 3070 688 3074 692
rect 3102 688 3106 692
rect 3358 688 3362 692
rect 3374 688 3378 692
rect 3398 688 3402 692
rect 3462 688 3466 692
rect 3494 688 3498 692
rect 3526 688 3530 692
rect 3590 688 3594 692
rect 3654 688 3658 692
rect 3710 688 3714 692
rect 86 678 90 682
rect 166 678 170 682
rect 206 678 210 682
rect 222 678 226 682
rect 238 678 242 682
rect 278 678 282 682
rect 318 678 322 682
rect 398 678 402 682
rect 414 678 418 682
rect 422 678 426 682
rect 486 678 490 682
rect 510 678 514 682
rect 734 678 738 682
rect 838 678 842 682
rect 974 678 978 682
rect 1150 678 1154 682
rect 1286 678 1290 682
rect 1350 678 1354 682
rect 1398 678 1402 682
rect 1478 678 1482 682
rect 1566 678 1570 682
rect 1742 678 1746 682
rect 1966 678 1970 682
rect 2118 678 2122 682
rect 2174 678 2178 682
rect 2622 678 2626 682
rect 2710 678 2714 682
rect 2726 678 2730 682
rect 2766 678 2770 682
rect 2822 678 2826 682
rect 2934 678 2938 682
rect 2950 678 2954 682
rect 3038 678 3042 682
rect 3262 678 3266 682
rect 3326 678 3330 682
rect 3366 678 3370 682
rect 3390 678 3394 682
rect 3430 678 3434 682
rect 3502 678 3506 682
rect 3534 678 3538 682
rect 3598 678 3602 682
rect 3606 678 3610 682
rect 3726 678 3730 682
rect 70 668 74 672
rect 198 668 202 672
rect 246 668 250 672
rect 262 668 266 672
rect 326 668 330 672
rect 438 668 442 672
rect 478 668 482 672
rect 526 668 530 672
rect 126 658 130 662
rect 182 658 186 662
rect 198 658 202 662
rect 254 658 258 662
rect 310 658 314 662
rect 374 658 378 662
rect 398 658 402 662
rect 446 658 450 662
rect 470 658 474 662
rect 518 658 522 662
rect 582 668 586 672
rect 718 668 722 672
rect 958 668 962 672
rect 1014 668 1018 672
rect 1134 668 1138 672
rect 1254 668 1258 672
rect 1262 668 1266 672
rect 1302 668 1306 672
rect 1318 668 1322 672
rect 1334 668 1338 672
rect 1350 668 1354 672
rect 1374 668 1378 672
rect 1598 668 1602 672
rect 1630 668 1634 672
rect 1726 668 1730 672
rect 1854 668 1858 672
rect 1886 668 1890 672
rect 1934 668 1938 672
rect 1950 668 1954 672
rect 1974 668 1978 672
rect 2006 668 2010 672
rect 590 658 594 662
rect 646 658 650 662
rect 774 658 778 662
rect 870 658 874 662
rect 958 658 962 662
rect 2046 668 2050 672
rect 2078 668 2082 672
rect 2142 668 2146 672
rect 2158 668 2162 672
rect 2166 668 2170 672
rect 2182 668 2186 672
rect 2262 668 2266 672
rect 2278 668 2282 672
rect 2294 668 2298 672
rect 2334 668 2338 672
rect 2350 668 2354 672
rect 2398 668 2402 672
rect 2430 668 2434 672
rect 2446 668 2450 672
rect 2462 668 2466 672
rect 2494 668 2498 672
rect 2526 668 2530 672
rect 2638 668 2642 672
rect 2734 668 2738 672
rect 2750 668 2754 672
rect 2782 668 2786 672
rect 2790 668 2794 672
rect 2830 668 2834 672
rect 2846 668 2850 672
rect 2878 668 2882 672
rect 2910 668 2914 672
rect 2974 668 2978 672
rect 3006 668 3010 672
rect 3022 668 3026 672
rect 3078 668 3082 672
rect 3094 668 3098 672
rect 3110 668 3114 672
rect 3158 668 3162 672
rect 3214 668 3218 672
rect 3254 668 3258 672
rect 3294 668 3298 672
rect 3310 668 3314 672
rect 3334 668 3338 672
rect 3454 668 3458 672
rect 3486 668 3490 672
rect 3518 668 3522 672
rect 3542 668 3546 672
rect 3558 668 3562 672
rect 3582 668 3586 672
rect 3630 668 3634 672
rect 3638 668 3642 672
rect 3662 668 3666 672
rect 3694 668 3698 672
rect 3710 668 3714 672
rect 3742 668 3746 672
rect 3758 668 3762 672
rect 3774 668 3778 672
rect 1086 658 1090 662
rect 1246 658 1250 662
rect 1278 658 1282 662
rect 1310 658 1314 662
rect 1358 658 1362 662
rect 1414 658 1418 662
rect 1446 658 1450 662
rect 1454 658 1458 662
rect 1494 658 1498 662
rect 1518 658 1522 662
rect 1534 658 1538 662
rect 1566 658 1570 662
rect 1590 658 1594 662
rect 1606 658 1610 662
rect 1638 658 1642 662
rect 1782 658 1786 662
rect 1926 658 1930 662
rect 1942 658 1946 662
rect 1982 658 1986 662
rect 1998 658 2002 662
rect 2022 658 2026 662
rect 2038 658 2042 662
rect 2102 658 2106 662
rect 2134 658 2138 662
rect 2150 658 2154 662
rect 2254 658 2258 662
rect 2286 658 2290 662
rect 2302 658 2306 662
rect 2310 658 2314 662
rect 2342 658 2346 662
rect 2366 658 2370 662
rect 2430 658 2434 662
rect 2438 658 2442 662
rect 2470 658 2474 662
rect 2502 658 2506 662
rect 2678 658 2682 662
rect 2710 658 2714 662
rect 2750 658 2754 662
rect 2782 658 2786 662
rect 2854 658 2858 662
rect 2886 658 2890 662
rect 2950 658 2954 662
rect 2998 658 3002 662
rect 3014 658 3018 662
rect 3030 658 3034 662
rect 3062 658 3066 662
rect 3078 658 3082 662
rect 3118 658 3122 662
rect 3126 658 3130 662
rect 3166 658 3170 662
rect 3206 658 3210 662
rect 3222 658 3226 662
rect 3286 658 3290 662
rect 3342 658 3346 662
rect 3382 658 3386 662
rect 3406 658 3410 662
rect 3430 658 3434 662
rect 3446 658 3450 662
rect 3478 658 3482 662
rect 3510 658 3514 662
rect 3550 658 3554 662
rect 3574 658 3578 662
rect 3630 658 3634 662
rect 3750 658 3754 662
rect 14 648 18 652
rect 390 648 394 652
rect 462 648 466 652
rect 686 650 690 654
rect 886 648 890 652
rect 910 648 914 652
rect 1102 650 1106 654
rect 1230 648 1234 652
rect 1318 648 1322 652
rect 1502 648 1506 652
rect 1574 648 1578 652
rect 1654 648 1658 652
rect 1678 648 1682 652
rect 1854 648 1858 652
rect 1894 648 1898 652
rect 1998 648 2002 652
rect 2022 648 2026 652
rect 2054 648 2058 652
rect 2086 648 2090 652
rect 2134 648 2138 652
rect 2318 648 2322 652
rect 2326 648 2330 652
rect 2358 648 2362 652
rect 2406 648 2410 652
rect 2478 648 2482 652
rect 2670 650 2674 654
rect 2846 648 2850 652
rect 2894 648 2898 652
rect 2974 648 2978 652
rect 2990 648 2994 652
rect 3062 648 3066 652
rect 3190 648 3194 652
rect 3270 648 3274 652
rect 3286 648 3290 652
rect 3470 648 3474 652
rect 3566 648 3570 652
rect 3654 648 3658 652
rect 3678 648 3682 652
rect 3758 648 3762 652
rect 1358 638 1362 642
rect 2822 638 2826 642
rect 126 627 130 631
rect 1102 627 1106 631
rect 2670 627 2674 631
rect 430 618 434 622
rect 446 618 450 622
rect 630 618 634 622
rect 686 618 690 622
rect 814 618 818 622
rect 910 618 914 622
rect 1054 618 1058 622
rect 1430 618 1434 622
rect 1462 618 1466 622
rect 1486 618 1490 622
rect 1678 618 1682 622
rect 1822 618 1826 622
rect 2014 618 2018 622
rect 2238 618 2242 622
rect 2278 618 2282 622
rect 2742 618 2746 622
rect 2942 618 2946 622
rect 3054 618 3058 622
rect 3142 618 3146 622
rect 3182 618 3186 622
rect 3206 618 3210 622
rect 3238 618 3242 622
rect 3326 618 3330 622
rect 3606 618 3610 622
rect 346 603 350 607
rect 353 603 357 607
rect 1362 603 1366 607
rect 1369 603 1373 607
rect 2386 603 2390 607
rect 2393 603 2397 607
rect 3410 603 3414 607
rect 3417 603 3421 607
rect 166 588 170 592
rect 374 588 378 592
rect 398 588 402 592
rect 550 588 554 592
rect 854 588 858 592
rect 1286 588 1290 592
rect 1334 588 1338 592
rect 1574 588 1578 592
rect 1694 588 1698 592
rect 1854 588 1858 592
rect 2414 588 2418 592
rect 2526 588 2530 592
rect 2670 588 2674 592
rect 2758 588 2762 592
rect 3454 588 3458 592
rect 3534 588 3538 592
rect 3614 588 3618 592
rect 3646 588 3650 592
rect 3678 588 3682 592
rect 3750 588 3754 592
rect 70 578 74 582
rect 646 578 650 582
rect 3174 578 3178 582
rect 406 568 410 572
rect 2270 568 2274 572
rect 3622 568 3626 572
rect 3654 568 3658 572
rect 3734 568 3738 572
rect 14 558 18 562
rect 38 556 42 560
rect 206 558 210 562
rect 214 558 218 562
rect 246 558 250 562
rect 278 558 282 562
rect 366 558 370 562
rect 390 558 394 562
rect 510 558 514 562
rect 678 556 682 560
rect 854 558 858 562
rect 1014 558 1018 562
rect 1054 558 1058 562
rect 1126 558 1130 562
rect 1150 558 1154 562
rect 1198 558 1202 562
rect 1214 558 1218 562
rect 1350 558 1354 562
rect 1438 558 1442 562
rect 1502 558 1506 562
rect 1558 558 1562 562
rect 1566 558 1570 562
rect 1646 558 1650 562
rect 1654 558 1658 562
rect 1854 558 1858 562
rect 1910 558 1914 562
rect 70 548 74 552
rect 190 548 194 552
rect 230 548 234 552
rect 278 548 282 552
rect 286 548 290 552
rect 302 548 306 552
rect 310 548 314 552
rect 398 548 402 552
rect 422 548 426 552
rect 502 548 506 552
rect 526 548 530 552
rect 542 548 546 552
rect 646 548 650 552
rect 742 548 746 552
rect 854 548 858 552
rect 958 548 962 552
rect 999 548 1003 552
rect 1078 548 1082 552
rect 1158 548 1162 552
rect 1174 548 1178 552
rect 1246 548 1250 552
rect 1278 548 1282 552
rect 1302 548 1306 552
rect 1310 548 1314 552
rect 1318 548 1322 552
rect 1414 548 1418 552
rect 1486 548 1490 552
rect 1510 548 1514 552
rect 1534 548 1538 552
rect 1542 548 1546 552
rect 1590 548 1594 552
rect 70 538 74 542
rect 182 538 186 542
rect 238 538 242 542
rect 270 538 274 542
rect 358 538 362 542
rect 382 538 386 542
rect 422 538 426 542
rect 454 538 458 542
rect 518 538 522 542
rect 534 538 538 542
rect 646 538 650 542
rect 822 538 826 542
rect 902 538 906 542
rect 1030 538 1034 542
rect 1038 538 1042 542
rect 1110 538 1114 542
rect 1126 538 1130 542
rect 1166 538 1170 542
rect 1182 538 1186 542
rect 1214 538 1218 542
rect 1366 538 1370 542
rect 1454 538 1458 542
rect 1478 538 1482 542
rect 1670 548 1674 552
rect 1702 548 1706 552
rect 1750 548 1754 552
rect 1950 558 1954 562
rect 1982 558 1986 562
rect 2062 558 2066 562
rect 2126 558 2130 562
rect 2230 558 2234 562
rect 2414 558 2418 562
rect 2454 558 2458 562
rect 2670 558 2674 562
rect 2694 558 2698 562
rect 2710 558 2714 562
rect 2798 558 2802 562
rect 2822 558 2826 562
rect 2862 558 2866 562
rect 2942 558 2946 562
rect 3022 558 3026 562
rect 3086 558 3090 562
rect 3158 558 3162 562
rect 3214 558 3218 562
rect 3254 558 3258 562
rect 3310 558 3314 562
rect 1998 548 2002 552
rect 2014 548 2018 552
rect 2102 548 2106 552
rect 2110 548 2114 552
rect 2134 548 2138 552
rect 2166 548 2170 552
rect 2206 548 2210 552
rect 2238 548 2242 552
rect 2262 548 2266 552
rect 2406 548 2410 552
rect 2438 548 2442 552
rect 2470 548 2474 552
rect 2502 548 2506 552
rect 2654 548 2658 552
rect 2678 548 2682 552
rect 2710 548 2714 552
rect 2726 548 2730 552
rect 2782 548 2786 552
rect 2862 548 2866 552
rect 2878 548 2882 552
rect 2910 548 2914 552
rect 2966 548 2970 552
rect 3006 548 3010 552
rect 3030 548 3034 552
rect 3070 548 3074 552
rect 3118 548 3122 552
rect 3126 548 3130 552
rect 3174 548 3178 552
rect 3198 548 3202 552
rect 3214 548 3218 552
rect 3222 548 3226 552
rect 3270 548 3274 552
rect 3294 548 3298 552
rect 3342 548 3346 552
rect 3358 548 3362 552
rect 3382 558 3386 562
rect 3566 558 3570 562
rect 3598 558 3602 562
rect 3606 558 3610 562
rect 3638 558 3642 562
rect 3766 558 3770 562
rect 3398 548 3402 552
rect 3446 548 3450 552
rect 3470 548 3474 552
rect 3486 548 3490 552
rect 3510 548 3514 552
rect 3534 548 3538 552
rect 3550 548 3554 552
rect 3566 548 3570 552
rect 3582 548 3586 552
rect 3598 548 3602 552
rect 3614 548 3618 552
rect 3646 548 3650 552
rect 3686 548 3690 552
rect 3710 548 3714 552
rect 3718 548 3722 552
rect 3734 548 3738 552
rect 3742 548 3746 552
rect 1550 538 1554 542
rect 1582 538 1586 542
rect 1598 538 1602 542
rect 1614 538 1618 542
rect 1622 538 1626 542
rect 1630 538 1634 542
rect 1646 538 1650 542
rect 1686 538 1690 542
rect 1806 538 1810 542
rect 1886 538 1890 542
rect 1910 538 1914 542
rect 1942 538 1946 542
rect 1974 538 1978 542
rect 2006 538 2010 542
rect 2046 538 2050 542
rect 2062 538 2066 542
rect 2086 538 2090 542
rect 2118 538 2122 542
rect 2142 538 2146 542
rect 2198 538 2202 542
rect 2214 538 2218 542
rect 2230 538 2234 542
rect 2366 538 2370 542
rect 2478 538 2482 542
rect 2518 538 2522 542
rect 2622 538 2626 542
rect 2718 538 2722 542
rect 2766 538 2770 542
rect 2774 538 2778 542
rect 2790 538 2794 542
rect 2806 538 2810 542
rect 2822 538 2826 542
rect 2846 538 2850 542
rect 2886 538 2890 542
rect 2918 538 2922 542
rect 2966 538 2970 542
rect 2974 538 2978 542
rect 3006 538 3010 542
rect 3038 538 3042 542
rect 3054 538 3058 542
rect 3094 538 3098 542
rect 3142 538 3146 542
rect 3182 538 3186 542
rect 3190 538 3194 542
rect 3230 538 3234 542
rect 3278 538 3282 542
rect 3286 538 3290 542
rect 3334 538 3338 542
rect 3350 538 3354 542
rect 3406 538 3410 542
rect 3446 538 3450 542
rect 3510 538 3514 542
rect 3542 538 3546 542
rect 3574 538 3578 542
rect 3742 538 3746 542
rect 86 528 90 532
rect 334 528 338 532
rect 430 528 434 532
rect 478 528 482 532
rect 630 528 634 532
rect 918 528 922 532
rect 1070 528 1074 532
rect 1102 528 1106 532
rect 1222 528 1226 532
rect 1262 528 1266 532
rect 1390 528 1394 532
rect 1430 528 1434 532
rect 1462 528 1466 532
rect 1470 528 1474 532
rect 1510 528 1514 532
rect 1686 528 1690 532
rect 1790 528 1794 532
rect 2070 528 2074 532
rect 2158 528 2162 532
rect 2350 528 2354 532
rect 2606 528 2610 532
rect 2830 528 2834 532
rect 2862 528 2866 532
rect 3054 528 3058 532
rect 3086 528 3090 532
rect 3430 528 3434 532
rect 3462 528 3466 532
rect 3486 528 3490 532
rect 3494 528 3498 532
rect 3518 528 3522 532
rect 3670 528 3674 532
rect 3694 528 3698 532
rect 3718 528 3722 532
rect 206 518 210 522
rect 214 518 218 522
rect 246 518 250 522
rect 494 518 498 522
rect 726 518 730 522
rect 758 518 762 522
rect 1022 518 1026 522
rect 1054 518 1058 522
rect 1094 518 1098 522
rect 1118 518 1122 522
rect 1150 518 1154 522
rect 1358 518 1362 522
rect 1398 518 1402 522
rect 1438 518 1442 522
rect 1598 518 1602 522
rect 1654 518 1658 522
rect 2030 518 2034 522
rect 2054 518 2058 522
rect 2150 518 2154 522
rect 2182 518 2186 522
rect 2486 518 2490 522
rect 2742 518 2746 522
rect 2814 518 2818 522
rect 2926 518 2930 522
rect 3022 518 3026 522
rect 3046 518 3050 522
rect 3238 518 3242 522
rect 3326 518 3330 522
rect 3374 518 3378 522
rect 850 503 854 507
rect 857 503 861 507
rect 1882 503 1886 507
rect 1889 503 1893 507
rect 2906 503 2910 507
rect 2913 503 2917 507
rect 166 488 170 492
rect 198 488 202 492
rect 238 488 242 492
rect 366 488 370 492
rect 406 488 410 492
rect 766 488 770 492
rect 1078 488 1082 492
rect 1102 488 1106 492
rect 1446 488 1450 492
rect 1686 488 1690 492
rect 1726 488 1730 492
rect 1750 488 1754 492
rect 1782 488 1786 492
rect 2390 488 2394 492
rect 2478 488 2482 492
rect 2558 488 2562 492
rect 2614 488 2618 492
rect 2830 488 2834 492
rect 3262 488 3266 492
rect 3542 488 3546 492
rect 3566 488 3570 492
rect 3630 488 3634 492
rect 3718 488 3722 492
rect 3742 488 3746 492
rect 86 478 90 482
rect 478 478 482 482
rect 670 478 674 482
rect 862 478 866 482
rect 998 478 1002 482
rect 1174 478 1178 482
rect 1366 478 1370 482
rect 1606 478 1610 482
rect 1710 478 1714 482
rect 1790 478 1794 482
rect 1830 478 1834 482
rect 1982 478 1986 482
rect 2070 478 2074 482
rect 2190 478 2194 482
rect 2310 478 2314 482
rect 2454 478 2458 482
rect 3134 478 3138 482
rect 3462 478 3466 482
rect 3558 478 3562 482
rect 3582 478 3586 482
rect 3598 478 3602 482
rect 3670 478 3674 482
rect 3726 478 3730 482
rect 3766 478 3770 482
rect 70 468 74 472
rect 182 468 186 472
rect 230 468 234 472
rect 294 468 298 472
rect 318 468 322 472
rect 342 468 346 472
rect 390 468 394 472
rect 446 468 450 472
rect 486 468 490 472
rect 518 468 522 472
rect 550 468 554 472
rect 686 468 690 472
rect 846 468 850 472
rect 982 468 986 472
rect 1094 468 1098 472
rect 1126 468 1130 472
rect 1134 468 1138 472
rect 1142 468 1146 472
rect 1198 468 1202 472
rect 1326 468 1330 472
rect 1342 468 1346 472
rect 1382 468 1386 472
rect 1414 468 1418 472
rect 1430 468 1434 472
rect 1438 468 1442 472
rect 1454 468 1458 472
rect 1518 468 1522 472
rect 1590 468 1594 472
rect 1718 468 1722 472
rect 1734 468 1738 472
rect 1758 468 1762 472
rect 1814 468 1818 472
rect 1830 468 1834 472
rect 1838 468 1842 472
rect 1854 468 1858 472
rect 1886 468 1890 472
rect 1918 468 1922 472
rect 1950 468 1954 472
rect 2086 468 2090 472
rect 2158 468 2162 472
rect 2206 468 2210 472
rect 2246 468 2250 472
rect 2278 468 2282 472
rect 2294 468 2298 472
rect 2310 468 2314 472
rect 2334 468 2338 472
rect 2374 468 2378 472
rect 2382 468 2386 472
rect 2414 468 2418 472
rect 2446 468 2450 472
rect 2462 468 2466 472
rect 2486 468 2490 472
rect 2502 468 2506 472
rect 2574 468 2578 472
rect 2598 468 2602 472
rect 2614 468 2618 472
rect 2654 468 2658 472
rect 2662 468 2666 472
rect 2718 468 2722 472
rect 2750 468 2754 472
rect 2782 468 2786 472
rect 2814 468 2818 472
rect 2822 468 2826 472
rect 2838 468 2842 472
rect 2870 468 2874 472
rect 2942 468 2946 472
rect 2974 468 2978 472
rect 2982 468 2986 472
rect 3038 468 3042 472
rect 3150 468 3154 472
rect 126 458 130 462
rect 254 458 258 462
rect 286 458 290 462
rect 294 458 298 462
rect 326 458 330 462
rect 382 458 386 462
rect 414 458 418 462
rect 422 458 426 462
rect 438 458 442 462
rect 462 458 466 462
rect 494 458 498 462
rect 518 458 522 462
rect 558 458 562 462
rect 726 458 730 462
rect 782 458 786 462
rect 806 458 810 462
rect 822 458 826 462
rect 894 458 898 462
rect 902 458 906 462
rect 950 458 954 462
rect 1038 458 1042 462
rect 1118 458 1122 462
rect 1150 458 1154 462
rect 1158 458 1162 462
rect 1166 458 1170 462
rect 1190 458 1194 462
rect 1206 458 1210 462
rect 1238 458 1242 462
rect 1246 458 1250 462
rect 1270 458 1274 462
rect 1286 458 1290 462
rect 1310 458 1314 462
rect 1350 458 1354 462
rect 1390 458 1394 462
rect 1422 458 1426 462
rect 1462 458 1466 462
rect 1486 458 1490 462
rect 1550 458 1554 462
rect 1646 458 1650 462
rect 1806 458 1810 462
rect 1846 458 1850 462
rect 1894 458 1898 462
rect 2030 458 2034 462
rect 2166 458 2170 462
rect 2214 458 2218 462
rect 2270 458 2274 462
rect 2286 458 2290 462
rect 2326 458 2330 462
rect 2366 458 2370 462
rect 2414 458 2418 462
rect 2438 458 2442 462
rect 2462 458 2466 462
rect 2494 458 2498 462
rect 2590 458 2594 462
rect 2622 458 2626 462
rect 2646 458 2650 462
rect 2654 458 2658 462
rect 2710 458 2714 462
rect 2742 458 2746 462
rect 2758 458 2762 462
rect 2814 458 2818 462
rect 2838 458 2842 462
rect 2854 458 2858 462
rect 2878 458 2882 462
rect 2934 458 2938 462
rect 2966 458 2970 462
rect 2990 458 2994 462
rect 3030 458 3034 462
rect 3150 458 3154 462
rect 3222 458 3226 462
rect 3238 458 3242 462
rect 3254 468 3258 472
rect 3270 468 3274 472
rect 3302 468 3306 472
rect 3358 468 3362 472
rect 3446 468 3450 472
rect 3606 468 3610 472
rect 3638 468 3642 472
rect 3654 468 3658 472
rect 3278 458 3282 462
rect 3350 458 3354 462
rect 3502 458 3506 462
rect 3574 458 3578 462
rect 3598 458 3602 462
rect 3614 458 3618 462
rect 3646 458 3650 462
rect 3686 458 3690 462
rect 3702 458 3706 462
rect 3734 458 3738 462
rect 38 450 42 454
rect 270 448 274 452
rect 302 448 306 452
rect 326 448 330 452
rect 398 448 402 452
rect 454 448 458 452
rect 510 448 514 452
rect 542 448 546 452
rect 574 448 578 452
rect 734 448 738 452
rect 814 448 818 452
rect 910 448 914 452
rect 934 448 938 452
rect 1278 448 1282 452
rect 1502 448 1506 452
rect 1542 448 1546 452
rect 1750 448 1754 452
rect 1782 448 1786 452
rect 1862 448 1866 452
rect 1910 448 1914 452
rect 1942 448 1946 452
rect 1974 448 1978 452
rect 2118 450 2122 454
rect 2222 448 2226 452
rect 2254 448 2258 452
rect 2342 448 2346 452
rect 2350 448 2354 452
rect 2438 448 2442 452
rect 2630 448 2634 452
rect 2686 448 2690 452
rect 2694 448 2698 452
rect 2710 448 2714 452
rect 2726 448 2730 452
rect 2790 448 2794 452
rect 2806 448 2810 452
rect 2862 448 2866 452
rect 2894 448 2898 452
rect 2950 448 2954 452
rect 2966 448 2970 452
rect 3014 448 3018 452
rect 3054 448 3058 452
rect 3182 450 3186 454
rect 3222 448 3226 452
rect 3294 448 3298 452
rect 3334 448 3338 452
rect 3398 448 3402 452
rect 3630 448 3634 452
rect 3662 448 3666 452
rect 526 438 530 442
rect 590 438 594 442
rect 798 438 802 442
rect 1110 438 1114 442
rect 1262 438 1266 442
rect 1342 438 1346 442
rect 1382 438 1386 442
rect 1414 438 1418 442
rect 1478 438 1482 442
rect 1486 438 1490 442
rect 126 427 130 431
rect 2646 428 2650 432
rect 3182 427 3186 431
rect 494 418 498 422
rect 558 418 562 422
rect 734 418 738 422
rect 934 418 938 422
rect 1254 418 1258 422
rect 1470 418 1474 422
rect 1542 418 1546 422
rect 1702 418 1706 422
rect 1798 418 1802 422
rect 1990 418 1994 422
rect 2118 418 2122 422
rect 2166 418 2170 422
rect 2238 418 2242 422
rect 2310 418 2314 422
rect 2366 418 2370 422
rect 2558 418 2562 422
rect 2582 418 2586 422
rect 2670 418 2674 422
rect 2742 418 2746 422
rect 2934 418 2938 422
rect 2990 418 2994 422
rect 3310 418 3314 422
rect 3398 418 3402 422
rect 346 403 350 407
rect 353 403 357 407
rect 1362 403 1366 407
rect 1369 403 1373 407
rect 2386 403 2390 407
rect 2393 403 2397 407
rect 3410 403 3414 407
rect 3417 403 3421 407
rect 14 388 18 392
rect 238 388 242 392
rect 262 388 266 392
rect 454 388 458 392
rect 486 388 490 392
rect 798 388 802 392
rect 1302 388 1306 392
rect 1454 388 1458 392
rect 1678 388 1682 392
rect 1822 388 1826 392
rect 1942 388 1946 392
rect 1966 388 1970 392
rect 2230 388 2234 392
rect 2422 388 2426 392
rect 2654 388 2658 392
rect 2894 388 2898 392
rect 2966 388 2970 392
rect 3110 388 3114 392
rect 3510 388 3514 392
rect 3534 388 3538 392
rect 3614 388 3618 392
rect 3630 388 3634 392
rect 3678 388 3682 392
rect 3726 388 3730 392
rect 142 378 146 382
rect 358 378 362 382
rect 926 378 930 382
rect 934 368 938 372
rect 966 368 970 372
rect 1030 368 1034 372
rect 1078 368 1082 372
rect 1142 368 1146 372
rect 1166 368 1170 372
rect 1870 368 1874 372
rect 2030 368 2034 372
rect 2086 368 2090 372
rect 2510 368 2514 372
rect 2758 368 2762 372
rect 3350 368 3354 372
rect 94 358 98 362
rect 310 358 314 362
rect 486 358 490 362
rect 798 358 802 362
rect 862 358 866 362
rect 910 358 914 362
rect 918 358 922 362
rect 1014 358 1018 362
rect 1046 358 1050 362
rect 1062 358 1066 362
rect 142 348 146 352
rect 358 348 362 352
rect 502 348 506 352
rect 590 348 594 352
rect 653 348 657 352
rect 750 348 754 352
rect 790 348 794 352
rect 846 348 850 352
rect 862 348 866 352
rect 870 348 874 352
rect 894 348 898 352
rect 926 348 930 352
rect 950 348 954 352
rect 990 348 994 352
rect 1022 348 1026 352
rect 1070 348 1074 352
rect 1094 348 1098 352
rect 1110 348 1114 352
rect 1134 348 1138 352
rect 1142 348 1146 352
rect 1198 358 1202 362
rect 1486 358 1490 362
rect 1526 358 1530 362
rect 1550 358 1554 362
rect 1574 358 1578 362
rect 1654 358 1658 362
rect 1678 358 1682 362
rect 1838 358 1842 362
rect 1854 358 1858 362
rect 1894 358 1898 362
rect 1974 358 1978 362
rect 2102 358 2106 362
rect 2198 358 2202 362
rect 2246 358 2250 362
rect 2310 358 2314 362
rect 2342 358 2346 362
rect 2374 358 2378 362
rect 2438 358 2442 362
rect 2454 358 2458 362
rect 2654 358 2658 362
rect 2710 358 2714 362
rect 2742 358 2746 362
rect 2814 358 2818 362
rect 1222 348 1226 352
rect 1278 348 1282 352
rect 1318 348 1322 352
rect 1350 348 1354 352
rect 1398 348 1402 352
rect 1406 348 1410 352
rect 1430 348 1434 352
rect 1446 348 1450 352
rect 1470 348 1474 352
rect 1478 348 1482 352
rect 1606 348 1610 352
rect 1638 348 1642 352
rect 1686 348 1690 352
rect 1870 348 1874 352
rect 1886 348 1890 352
rect 1982 348 1986 352
rect 2014 348 2018 352
rect 2022 348 2026 352
rect 2062 348 2066 352
rect 2078 348 2082 352
rect 2126 348 2130 352
rect 2190 348 2194 352
rect 2214 348 2218 352
rect 2262 348 2266 352
rect 2302 348 2306 352
rect 2334 348 2338 352
rect 2390 348 2394 352
rect 2398 348 2402 352
rect 2462 348 2466 352
rect 2494 348 2498 352
rect 2638 348 2642 352
rect 2654 348 2658 352
rect 2702 348 2706 352
rect 2726 348 2730 352
rect 2758 348 2762 352
rect 2766 348 2770 352
rect 2798 348 2802 352
rect 2854 358 2858 362
rect 2942 358 2946 362
rect 2966 358 2970 362
rect 3158 358 3162 362
rect 3214 358 3218 362
rect 2878 348 2882 352
rect 2926 348 2930 352
rect 2974 348 2978 352
rect 3126 348 3130 352
rect 3174 348 3178 352
rect 3198 348 3202 352
rect 3254 358 3258 362
rect 3302 358 3306 362
rect 3334 358 3338 362
rect 3366 358 3370 362
rect 3470 358 3474 362
rect 3502 358 3506 362
rect 3638 358 3642 362
rect 3270 348 3274 352
rect 3318 348 3322 352
rect 3350 348 3354 352
rect 3382 348 3386 352
rect 3390 348 3394 352
rect 3446 348 3450 352
rect 3470 348 3474 352
rect 3486 348 3490 352
rect 3622 348 3626 352
rect 3646 348 3650 352
rect 3654 348 3658 352
rect 3662 348 3666 352
rect 70 338 74 342
rect 142 338 146 342
rect 358 338 362 342
rect 534 338 538 342
rect 750 338 754 342
rect 838 338 842 342
rect 878 338 882 342
rect 910 338 914 342
rect 982 338 986 342
rect 998 338 1002 342
rect 1102 338 1106 342
rect 1118 338 1122 342
rect 1134 338 1138 342
rect 1190 338 1194 342
rect 1246 338 1250 342
rect 1326 338 1330 342
rect 1390 338 1394 342
rect 1502 338 1506 342
rect 1510 338 1514 342
rect 1534 338 1538 342
rect 1558 338 1562 342
rect 1598 338 1602 342
rect 1654 338 1658 342
rect 1726 338 1730 342
rect 1838 338 1842 342
rect 1862 338 1866 342
rect 1950 338 1954 342
rect 1990 338 1994 342
rect 2006 338 2010 342
rect 2022 338 2026 342
rect 2046 338 2050 342
rect 2086 338 2090 342
rect 2166 338 2170 342
rect 2238 338 2242 342
rect 2254 338 2258 342
rect 2270 338 2274 342
rect 2286 338 2290 342
rect 2294 338 2298 342
rect 2334 338 2338 342
rect 2350 338 2354 342
rect 2366 338 2370 342
rect 2414 338 2418 342
rect 2430 338 2434 342
rect 2470 338 2474 342
rect 2502 338 2506 342
rect 2606 338 2610 342
rect 2694 338 2698 342
rect 2718 338 2722 342
rect 2734 338 2738 342
rect 2766 338 2770 342
rect 2774 338 2778 342
rect 2790 338 2794 342
rect 2822 338 2826 342
rect 2878 338 2882 342
rect 2886 338 2890 342
rect 2910 338 2914 342
rect 2934 338 2938 342
rect 3014 338 3018 342
rect 3134 338 3138 342
rect 3166 338 3170 342
rect 3182 338 3186 342
rect 3190 338 3194 342
rect 3222 338 3226 342
rect 3278 338 3282 342
rect 3286 338 3290 342
rect 3326 338 3330 342
rect 3374 338 3378 342
rect 3390 338 3394 342
rect 3406 338 3410 342
rect 3422 338 3426 342
rect 3438 338 3442 342
rect 3478 338 3482 342
rect 3518 338 3522 342
rect 3590 338 3594 342
rect 3670 338 3674 342
rect 3710 338 3714 342
rect 3758 338 3762 342
rect 158 328 162 332
rect 286 328 290 332
rect 374 328 378 332
rect 550 328 554 332
rect 734 328 738 332
rect 822 328 826 332
rect 1046 328 1050 332
rect 1374 328 1378 332
rect 1422 328 1426 332
rect 1590 328 1594 332
rect 1622 328 1626 332
rect 1742 328 1746 332
rect 1926 328 1930 332
rect 2062 328 2066 332
rect 2110 328 2114 332
rect 2142 328 2146 332
rect 2166 328 2170 332
rect 2278 328 2282 332
rect 2310 328 2314 332
rect 2470 328 2474 332
rect 2590 328 2594 332
rect 2678 328 2682 332
rect 3030 328 3034 332
rect 3150 328 3154 332
rect 3294 328 3298 332
rect 3302 328 3306 332
rect 3422 328 3426 332
rect 3598 328 3602 332
rect 3622 328 3626 332
rect 630 318 634 322
rect 966 318 970 322
rect 1078 318 1082 322
rect 1238 318 1242 322
rect 1302 318 1306 322
rect 1334 318 1338 322
rect 1494 318 1498 322
rect 1526 318 1530 322
rect 1550 318 1554 322
rect 1574 318 1578 322
rect 1998 318 2002 322
rect 2070 318 2074 322
rect 2478 318 2482 322
rect 2686 318 2690 322
rect 2846 318 2850 322
rect 3142 318 3146 322
rect 3246 318 3250 322
rect 3502 318 3506 322
rect 850 303 854 307
rect 857 303 861 307
rect 1882 303 1886 307
rect 1889 303 1893 307
rect 2906 303 2910 307
rect 2913 303 2917 307
rect 166 288 170 292
rect 638 288 642 292
rect 1046 288 1050 292
rect 1214 288 1218 292
rect 1398 288 1402 292
rect 1446 288 1450 292
rect 1862 288 1866 292
rect 1934 288 1938 292
rect 2022 288 2026 292
rect 2046 288 2050 292
rect 2294 288 2298 292
rect 2342 288 2346 292
rect 2510 288 2514 292
rect 2550 288 2554 292
rect 2622 288 2626 292
rect 2822 288 2826 292
rect 3110 288 3114 292
rect 3590 288 3594 292
rect 3614 288 3618 292
rect 86 278 90 282
rect 270 278 274 282
rect 462 278 466 282
rect 830 278 834 282
rect 974 278 978 282
rect 1134 278 1138 282
rect 1318 278 1322 282
rect 1966 278 1970 282
rect 2078 278 2082 282
rect 2118 278 2122 282
rect 2150 278 2154 282
rect 2214 278 2218 282
rect 2422 278 2426 282
rect 2614 278 2618 282
rect 2718 278 2722 282
rect 2942 278 2946 282
rect 2982 278 2986 282
rect 3190 278 3194 282
rect 3334 278 3338 282
rect 3342 278 3346 282
rect 3446 278 3450 282
rect 3694 278 3698 282
rect 70 268 74 272
rect 286 268 290 272
rect 422 268 426 272
rect 478 268 482 272
rect 550 268 554 272
rect 582 268 586 272
rect 678 268 682 272
rect 749 268 753 272
rect 846 268 850 272
rect 934 268 938 272
rect 950 268 954 272
rect 1014 268 1018 272
rect 1062 268 1066 272
rect 1070 268 1074 272
rect 1166 268 1170 272
rect 1182 268 1186 272
rect 1302 268 1306 272
rect 1518 268 1522 272
rect 1534 268 1538 272
rect 1590 268 1594 272
rect 1614 268 1618 272
rect 1662 268 1666 272
rect 1678 268 1682 272
rect 1734 268 1738 272
rect 1750 268 1754 272
rect 1806 268 1810 272
rect 1822 268 1826 272
rect 1838 268 1842 272
rect 1878 268 1882 272
rect 1902 268 1906 272
rect 1926 268 1930 272
rect 1958 268 1962 272
rect 1974 268 1978 272
rect 1990 268 1994 272
rect 2030 268 2034 272
rect 2038 268 2042 272
rect 2062 268 2066 272
rect 2110 268 2114 272
rect 2134 268 2138 272
rect 2206 268 2210 272
rect 2238 268 2242 272
rect 2246 268 2250 272
rect 2286 268 2290 272
rect 2302 268 2306 272
rect 2438 268 2442 272
rect 2526 268 2530 272
rect 2542 268 2546 272
rect 2558 268 2562 272
rect 2582 268 2586 272
rect 2598 268 2602 272
rect 2702 268 2706 272
rect 2854 268 2858 272
rect 2862 268 2866 272
rect 2910 268 2914 272
rect 2942 268 2946 272
rect 2958 268 2962 272
rect 2974 268 2978 272
rect 3014 268 3018 272
rect 126 258 130 262
rect 334 258 338 262
rect 518 258 522 262
rect 558 258 562 262
rect 694 258 698 262
rect 790 258 794 262
rect 846 258 850 262
rect 942 258 946 262
rect 958 258 962 262
rect 990 258 994 262
rect 1022 258 1026 262
rect 1078 258 1082 262
rect 1110 258 1114 262
rect 1150 258 1154 262
rect 1158 258 1162 262
rect 1230 258 1234 262
rect 1254 258 1258 262
rect 1358 258 1362 262
rect 1438 258 1442 262
rect 1462 258 1466 262
rect 1470 258 1474 262
rect 1494 258 1498 262
rect 1510 258 1514 262
rect 1542 258 1546 262
rect 1566 258 1570 262
rect 1582 258 1586 262
rect 1614 258 1618 262
rect 1630 258 1634 262
rect 1654 258 1658 262
rect 1670 258 1674 262
rect 1686 258 1690 262
rect 1702 258 1706 262
rect 1726 258 1730 262
rect 1742 258 1746 262
rect 1758 258 1762 262
rect 1774 258 1778 262
rect 1798 258 1802 262
rect 1814 258 1818 262
rect 1830 258 1834 262
rect 1950 258 1954 262
rect 1982 258 1986 262
rect 2102 258 2106 262
rect 2126 258 2130 262
rect 2182 258 2186 262
rect 2198 258 2202 262
rect 2230 258 2234 262
rect 2254 258 2258 262
rect 2278 258 2282 262
rect 2310 258 2314 262
rect 2382 258 2386 262
rect 2486 258 2490 262
rect 2534 258 2538 262
rect 2566 258 2570 262
rect 2574 258 2578 262
rect 2590 258 2594 262
rect 2606 258 2610 262
rect 2630 258 2634 262
rect 2654 258 2658 262
rect 2799 258 2803 262
rect 2846 258 2850 262
rect 2870 258 2874 262
rect 2926 258 2930 262
rect 3006 258 3010 262
rect 3022 258 3026 262
rect 3038 258 3042 262
rect 3054 268 3058 272
rect 3070 268 3074 272
rect 3206 268 3210 272
rect 3278 268 3282 272
rect 3318 268 3322 272
rect 3462 268 3466 272
rect 3534 268 3538 272
rect 3710 268 3714 272
rect 3078 258 3082 262
rect 3150 258 3154 262
rect 3286 258 3290 262
rect 3310 258 3314 262
rect 3326 258 3330 262
rect 3462 258 3466 262
rect 3494 258 3498 262
rect 3710 258 3714 262
rect 38 250 42 254
rect 318 250 322 254
rect 510 250 514 254
rect 574 248 578 252
rect 654 248 658 252
rect 710 248 714 252
rect 894 248 898 252
rect 958 248 962 252
rect 982 248 986 252
rect 1038 248 1042 252
rect 1046 248 1050 252
rect 1102 248 1106 252
rect 1174 248 1178 252
rect 1198 248 1202 252
rect 1254 248 1258 252
rect 1502 248 1506 252
rect 1574 248 1578 252
rect 1590 248 1594 252
rect 1622 248 1626 252
rect 1694 248 1698 252
rect 1766 248 1770 252
rect 1942 248 1946 252
rect 2006 248 2010 252
rect 2014 248 2018 252
rect 2102 248 2106 252
rect 2182 248 2186 252
rect 2214 248 2218 252
rect 2270 248 2274 252
rect 2470 250 2474 254
rect 2510 248 2514 252
rect 2670 250 2674 254
rect 2830 248 2834 252
rect 2846 248 2850 252
rect 2886 248 2890 252
rect 2894 248 2898 252
rect 2990 248 2994 252
rect 3022 248 3026 252
rect 3094 248 3098 252
rect 3254 248 3258 252
rect 3302 248 3306 252
rect 3510 248 3514 252
rect 3742 250 3746 254
rect 998 238 1002 242
rect 1022 238 1026 242
rect 1118 238 1122 242
rect 1182 238 1186 242
rect 1486 238 1490 242
rect 1534 238 1538 242
rect 1558 238 1562 242
rect 1638 238 1642 242
rect 1710 238 1714 242
rect 1782 238 1786 242
rect 1862 238 1866 242
rect 1886 238 1890 242
rect 1926 238 1930 242
rect 1990 238 1994 242
rect 2942 238 2946 242
rect 126 227 130 231
rect 2470 227 2474 231
rect 2670 227 2674 231
rect 3742 227 3746 231
rect 190 218 194 222
rect 318 218 322 222
rect 382 218 386 222
rect 510 218 514 222
rect 558 218 562 222
rect 638 218 642 222
rect 670 218 674 222
rect 734 218 738 222
rect 894 218 898 222
rect 990 218 994 222
rect 1078 218 1082 222
rect 1254 218 1258 222
rect 1478 218 1482 222
rect 1566 218 1570 222
rect 1630 218 1634 222
rect 1702 218 1706 222
rect 1774 218 1778 222
rect 1846 218 1850 222
rect 2254 218 2258 222
rect 2870 218 2874 222
rect 3006 218 3010 222
rect 3062 218 3066 222
rect 3078 218 3082 222
rect 3254 218 3258 222
rect 3286 218 3290 222
rect 3510 218 3514 222
rect 3590 218 3594 222
rect 346 203 350 207
rect 353 203 357 207
rect 1362 203 1366 207
rect 1369 203 1373 207
rect 2386 203 2390 207
rect 2393 203 2397 207
rect 3410 203 3414 207
rect 3417 203 3421 207
rect 86 188 90 192
rect 110 188 114 192
rect 446 188 450 192
rect 590 188 594 192
rect 1318 188 1322 192
rect 1462 188 1466 192
rect 1630 188 1634 192
rect 2078 188 2082 192
rect 2198 188 2202 192
rect 2438 188 2442 192
rect 2478 188 2482 192
rect 2622 188 2626 192
rect 2742 188 2746 192
rect 2854 188 2858 192
rect 3062 188 3066 192
rect 3206 188 3210 192
rect 3302 188 3306 192
rect 3470 188 3474 192
rect 3518 188 3522 192
rect 3582 188 3586 192
rect 3646 188 3650 192
rect 3718 188 3722 192
rect 3742 188 3746 192
rect 934 179 938 183
rect 1030 178 1034 182
rect 1038 168 1042 172
rect 1094 168 1098 172
rect 1270 178 1274 182
rect 1790 179 1794 183
rect 1950 179 1954 183
rect 2310 179 2314 183
rect 1134 168 1138 172
rect 1654 168 1658 172
rect 2830 168 2834 172
rect 3550 168 3554 172
rect 3710 168 3714 172
rect 446 158 450 162
rect 614 158 618 162
rect 630 158 634 162
rect 662 158 666 162
rect 718 158 722 162
rect 750 158 754 162
rect 934 156 938 160
rect 982 158 986 162
rect 998 158 1002 162
rect 1022 158 1026 162
rect 1062 158 1066 162
rect 1078 158 1082 162
rect 1110 158 1114 162
rect 1190 158 1194 162
rect 1318 158 1322 162
rect 1630 158 1634 162
rect 1790 156 1794 160
rect 1814 158 1818 162
rect 22 148 26 152
rect 94 148 98 152
rect 190 148 194 152
rect 550 148 554 152
rect 598 148 602 152
rect 646 148 650 152
rect 702 148 706 152
rect 726 148 730 152
rect 846 148 850 152
rect 958 148 962 152
rect 982 148 986 152
rect 998 148 1002 152
rect 1030 148 1034 152
rect 1062 148 1066 152
rect 1102 148 1106 152
rect 1174 148 1178 152
rect 1190 148 1194 152
rect 1214 148 1218 152
rect 1246 148 1250 152
rect 1318 148 1322 152
rect 1526 148 1530 152
rect 1702 148 1706 152
rect 1950 156 1954 160
rect 2118 158 2122 162
rect 1934 148 1938 152
rect 2102 148 2106 152
rect 2182 158 2186 162
rect 2190 158 2194 162
rect 2206 158 2210 162
rect 2246 158 2250 162
rect 2310 156 2314 160
rect 2622 158 2626 162
rect 2702 158 2706 162
rect 2950 158 2954 162
rect 2958 158 2962 162
rect 3014 158 3018 162
rect 3206 158 3210 162
rect 3470 158 3474 162
rect 3566 158 3570 162
rect 3726 158 3730 162
rect 2142 148 2146 152
rect 2166 148 2170 152
rect 2182 148 2186 152
rect 2230 148 2234 152
rect 2262 148 2266 152
rect 2294 148 2298 152
rect 2398 148 2402 152
rect 2518 148 2522 152
rect 2630 148 2634 152
rect 2662 148 2666 152
rect 2718 148 2722 152
rect 2846 148 2850 152
rect 2878 148 2882 152
rect 2926 148 2930 152
rect 2934 148 2938 152
rect 2958 148 2962 152
rect 2974 148 2978 152
rect 2998 148 3002 152
rect 3014 148 3018 152
rect 3046 148 3050 152
rect 3190 148 3194 152
rect 3366 148 3370 152
rect 3462 148 3466 152
rect 3534 148 3538 152
rect 3558 148 3562 152
rect 3598 148 3602 152
rect 3630 148 3634 152
rect 3662 148 3666 152
rect 3670 148 3674 152
rect 3718 148 3722 152
rect 3758 148 3762 152
rect 6 138 10 142
rect 30 138 34 142
rect 166 138 170 142
rect 198 138 202 142
rect 270 138 274 142
rect 334 138 338 142
rect 342 138 346 142
rect 494 138 498 142
rect 606 138 610 142
rect 638 138 642 142
rect 694 138 698 142
rect 710 138 714 142
rect 726 138 730 142
rect 902 138 906 142
rect 974 138 978 142
rect 1014 138 1018 142
rect 1054 138 1058 142
rect 1142 138 1146 142
rect 1198 138 1202 142
rect 1222 138 1226 142
rect 1366 138 1370 142
rect 1422 138 1426 142
rect 1582 138 1586 142
rect 1758 138 1762 142
rect 1830 138 1834 142
rect 1894 138 1898 142
rect 1982 138 1986 142
rect 2094 138 2098 142
rect 2150 138 2154 142
rect 2158 138 2162 142
rect 2206 138 2210 142
rect 2238 138 2242 142
rect 2254 138 2258 142
rect 2270 138 2274 142
rect 2342 138 2346 142
rect 2574 138 2578 142
rect 2686 138 2690 142
rect 2726 138 2730 142
rect 2798 138 2802 142
rect 2838 138 2842 142
rect 2982 138 2986 142
rect 2990 138 2994 142
rect 3030 138 3034 142
rect 3038 138 3042 142
rect 3158 138 3162 142
rect 3230 138 3234 142
rect 3294 138 3298 142
rect 3310 138 3314 142
rect 3422 138 3426 142
rect 3606 138 3610 142
rect 3678 138 3682 142
rect 30 128 34 132
rect 510 128 514 132
rect 806 128 810 132
rect 886 128 890 132
rect 1158 128 1162 132
rect 1206 128 1210 132
rect 1382 128 1386 132
rect 1566 128 1570 132
rect 1742 128 1746 132
rect 1998 128 2002 132
rect 2358 128 2362 132
rect 2558 128 2562 132
rect 2646 128 2650 132
rect 3022 128 3026 132
rect 3142 128 3146 132
rect 3406 128 3410 132
rect 3694 128 3698 132
rect 174 118 178 122
rect 254 118 258 122
rect 414 118 418 122
rect 686 118 690 122
rect 782 118 786 122
rect 1486 118 1490 122
rect 2126 118 2130 122
rect 2214 118 2218 122
rect 2678 118 2682 122
rect 2950 118 2954 122
rect 3550 118 3554 122
rect 3686 118 3690 122
rect 850 103 854 107
rect 857 103 861 107
rect 1882 103 1886 107
rect 1889 103 1893 107
rect 2906 103 2910 107
rect 2913 103 2917 107
rect 230 88 234 92
rect 278 88 282 92
rect 1462 88 1466 92
rect 2198 88 2202 92
rect 2374 88 2378 92
rect 2590 88 2594 92
rect 2838 88 2842 92
rect 3086 88 3090 92
rect 3110 88 3114 92
rect 3126 88 3130 92
rect 3150 88 3154 92
rect 3334 88 3338 92
rect 3430 88 3434 92
rect 3454 88 3458 92
rect 3502 88 3506 92
rect 3614 88 3618 92
rect 3638 88 3642 92
rect 3662 88 3666 92
rect 3718 88 3722 92
rect 118 78 122 82
rect 486 78 490 82
rect 734 78 738 82
rect 918 78 922 82
rect 1118 78 1122 82
rect 1318 78 1322 82
rect 1630 78 1634 82
rect 1918 78 1922 82
rect 2006 78 2010 82
rect 2094 78 2098 82
rect 2294 78 2298 82
rect 2494 78 2498 82
rect 2670 78 2674 82
rect 2854 78 2858 82
rect 2870 78 2874 82
rect 134 68 138 72
rect 182 58 186 62
rect 222 58 226 62
rect 502 68 506 72
rect 750 68 754 72
rect 902 68 906 72
rect 1102 68 1106 72
rect 1158 68 1162 72
rect 1302 68 1306 72
rect 1518 68 1522 72
rect 1614 68 1618 72
rect 1750 68 1754 72
rect 1814 68 1818 72
rect 1902 68 1906 72
rect 2078 68 2082 72
rect 2134 68 2138 72
rect 2175 68 2179 72
rect 2206 68 2210 72
rect 2278 68 2282 72
rect 2510 68 2514 72
rect 2630 68 2634 72
rect 2686 68 2690 72
rect 2758 68 2762 72
rect 2822 68 2826 72
rect 3006 78 3010 82
rect 3102 78 3106 82
rect 3134 78 3138 82
rect 3230 78 3234 82
rect 3606 78 3610 82
rect 3630 78 3634 82
rect 3726 78 3730 82
rect 2886 68 2890 72
rect 2894 68 2898 72
rect 2990 68 2994 72
rect 3246 68 3250 72
rect 3350 68 3354 72
rect 3526 68 3530 72
rect 3574 68 3578 72
rect 3582 68 3586 72
rect 3686 68 3690 72
rect 3702 68 3706 72
rect 3758 68 3762 72
rect 262 58 266 62
rect 302 58 306 62
rect 326 58 330 62
rect 350 58 354 62
rect 550 58 554 62
rect 590 58 594 62
rect 598 58 602 62
rect 622 58 626 62
rect 653 58 657 62
rect 790 58 794 62
rect 958 58 962 62
rect 1054 58 1058 62
rect 1254 58 1258 62
rect 1526 58 1530 62
rect 1566 58 1570 62
rect 1958 58 1962 62
rect 2038 58 2042 62
rect 2230 58 2234 62
rect 2558 58 2562 62
rect 2734 58 2738 62
rect 2830 58 2834 62
rect 2854 58 2858 62
rect 2902 58 2906 62
rect 3046 58 3050 62
rect 3118 58 3122 62
rect 3190 58 3194 62
rect 3302 58 3306 62
rect 3334 58 3338 62
rect 3390 58 3394 62
rect 3446 58 3450 62
rect 3470 58 3474 62
rect 3486 58 3490 62
rect 3542 58 3546 62
rect 3622 58 3626 62
rect 3646 58 3650 62
rect 3678 58 3682 62
rect 3694 58 3698 62
rect 3726 58 3730 62
rect 3750 58 3754 62
rect 182 48 186 52
rect 230 48 234 52
rect 254 48 258 52
rect 534 50 538 54
rect 798 48 802 52
rect 854 48 858 52
rect 1054 48 1058 52
rect 1254 48 1258 52
rect 1582 50 1586 54
rect 1870 50 1874 54
rect 2046 50 2050 54
rect 2190 48 2194 52
rect 2246 50 2250 54
rect 2414 48 2418 52
rect 2542 50 2546 54
rect 2734 48 2738 52
rect 2942 48 2946 52
rect 3294 48 3298 52
rect 3342 48 3346 52
rect 3350 48 3354 52
rect 3366 48 3370 52
rect 3398 48 3402 52
rect 3478 48 3482 52
rect 3710 48 3714 52
rect 3734 48 3738 52
rect 6 38 10 42
rect 270 38 274 42
rect 3326 38 3330 42
rect 3382 38 3386 42
rect 3462 38 3466 42
rect 534 27 538 31
rect 1582 27 1586 31
rect 1870 27 1874 31
rect 2542 27 2546 31
rect 3390 28 3394 32
rect 3590 28 3594 32
rect 182 18 186 22
rect 206 18 210 22
rect 286 18 290 22
rect 310 18 314 22
rect 334 18 338 22
rect 374 18 378 22
rect 574 18 578 22
rect 614 18 618 22
rect 638 18 642 22
rect 798 18 802 22
rect 854 18 858 22
rect 1030 18 1034 22
rect 1054 18 1058 22
rect 1230 18 1234 22
rect 1254 18 1258 22
rect 1446 18 1450 22
rect 1542 18 1546 22
rect 1742 18 1746 22
rect 2046 18 2050 22
rect 2246 18 2250 22
rect 2734 18 2738 22
rect 2942 18 2946 22
rect 3294 18 3298 22
rect 346 3 350 7
rect 353 3 357 7
rect 1362 3 1366 7
rect 1369 3 1373 7
rect 2386 3 2390 7
rect 2393 3 2397 7
rect 3410 3 3414 7
rect 3417 3 3421 7
<< metal2 >>
rect 158 3631 162 3632
rect 214 3631 218 3632
rect 150 3628 162 3631
rect 206 3628 218 3631
rect 254 3631 258 3632
rect 278 3631 282 3632
rect 302 3631 306 3632
rect 326 3631 330 3632
rect 254 3628 265 3631
rect 150 3592 153 3628
rect 66 3538 70 3541
rect 82 3538 86 3541
rect 6 3472 9 3538
rect 30 3472 33 3538
rect 102 3472 105 3538
rect 166 3531 169 3548
rect 174 3542 177 3548
rect 166 3528 177 3531
rect 6 3442 9 3448
rect 22 3402 25 3458
rect 134 3432 137 3518
rect 166 3472 169 3478
rect 86 3422 89 3428
rect 174 3412 177 3528
rect 206 3492 209 3628
rect 262 3592 265 3628
rect 270 3628 282 3631
rect 294 3628 306 3631
rect 318 3628 330 3631
rect 430 3628 434 3632
rect 542 3631 546 3632
rect 534 3628 546 3631
rect 742 3631 746 3632
rect 766 3631 770 3632
rect 742 3628 753 3631
rect 270 3592 273 3628
rect 294 3592 297 3628
rect 318 3592 321 3628
rect 344 3603 346 3607
rect 350 3603 353 3607
rect 357 3603 360 3607
rect 430 3602 433 3628
rect 534 3592 537 3628
rect 750 3592 753 3628
rect 758 3628 770 3631
rect 886 3628 890 3632
rect 958 3628 962 3632
rect 982 3631 986 3632
rect 982 3628 993 3631
rect 758 3592 761 3628
rect 886 3602 889 3628
rect 494 3560 497 3579
rect 694 3560 697 3579
rect 934 3560 937 3579
rect 314 3548 318 3551
rect 514 3548 518 3551
rect 730 3548 734 3551
rect 238 3532 241 3538
rect 198 3452 201 3458
rect 182 3392 185 3418
rect 6 3372 9 3378
rect 30 3362 33 3368
rect 222 3362 225 3388
rect 246 3372 249 3548
rect 286 3522 289 3548
rect 318 3472 321 3478
rect 334 3462 337 3468
rect 366 3431 369 3450
rect 294 3392 297 3408
rect 344 3403 346 3407
rect 350 3403 353 3407
rect 357 3403 360 3407
rect 326 3392 329 3398
rect 374 3392 377 3548
rect 446 3522 449 3528
rect 422 3492 425 3508
rect 382 3392 385 3458
rect 438 3452 441 3458
rect 454 3402 457 3418
rect 286 3352 289 3388
rect 6 3242 9 3248
rect 10 3138 14 3141
rect 6 3042 9 3048
rect 6 2942 9 2948
rect 14 2872 17 3138
rect 22 3082 25 3348
rect 54 3342 57 3348
rect 74 3338 77 3341
rect 54 3332 57 3338
rect 66 3328 70 3331
rect 158 3311 161 3328
rect 174 3322 177 3338
rect 206 3312 209 3348
rect 246 3342 249 3348
rect 254 3332 257 3348
rect 270 3332 273 3348
rect 310 3342 313 3358
rect 318 3352 321 3388
rect 346 3358 350 3361
rect 266 3318 270 3321
rect 278 3312 281 3338
rect 158 3308 169 3311
rect 118 3252 121 3278
rect 134 3262 137 3268
rect 134 3192 137 3248
rect 74 3138 78 3141
rect 42 3078 46 3081
rect 22 3052 25 3058
rect 22 2932 25 2948
rect 78 2942 81 3138
rect 166 3132 169 3308
rect 174 3262 177 3308
rect 286 3302 289 3338
rect 318 3302 321 3338
rect 222 3292 225 3298
rect 174 3152 177 3258
rect 182 3222 185 3248
rect 206 3242 209 3258
rect 206 3222 209 3238
rect 270 3231 273 3250
rect 302 3232 305 3268
rect 318 3252 321 3278
rect 358 3262 361 3388
rect 406 3382 409 3388
rect 370 3348 374 3351
rect 366 3302 369 3338
rect 374 3302 377 3348
rect 390 3332 393 3358
rect 366 3282 369 3298
rect 398 3292 401 3338
rect 414 3292 417 3318
rect 402 3288 406 3291
rect 358 3221 361 3258
rect 422 3242 425 3348
rect 442 3328 446 3331
rect 454 3292 457 3368
rect 446 3262 449 3268
rect 434 3248 438 3251
rect 358 3218 369 3221
rect 344 3203 346 3207
rect 350 3203 353 3207
rect 357 3203 360 3207
rect 182 3160 185 3179
rect 358 3162 361 3188
rect 118 3012 121 3078
rect 134 3062 137 3068
rect 86 2992 89 3008
rect 166 2952 169 3128
rect 174 3062 177 3148
rect 214 3142 217 3158
rect 366 3152 369 3218
rect 454 3212 457 3248
rect 274 3148 278 3151
rect 230 3122 233 3128
rect 206 3072 209 3078
rect 230 3072 233 3078
rect 218 3068 222 3071
rect 238 3062 241 3068
rect 226 3058 230 3061
rect 254 3052 257 3098
rect 242 3048 246 3051
rect 182 3022 185 3048
rect 230 2992 233 3038
rect 98 2938 102 2941
rect 170 2938 174 2941
rect 242 2938 246 2941
rect 30 2912 33 2938
rect 30 2882 33 2888
rect 54 2872 57 2878
rect 6 2842 9 2848
rect 6 2742 9 2748
rect 6 2662 9 2668
rect 6 2562 9 2568
rect 6 2482 9 2488
rect 6 2452 9 2468
rect 6 2342 9 2348
rect 14 2272 17 2868
rect 26 2858 30 2861
rect 58 2858 62 2861
rect 46 2852 49 2858
rect 62 2842 65 2848
rect 70 2822 73 2908
rect 54 2482 57 2798
rect 70 2672 73 2818
rect 78 2712 81 2848
rect 86 2812 89 2918
rect 94 2882 97 2888
rect 118 2872 121 2878
rect 122 2858 126 2861
rect 110 2852 113 2858
rect 130 2848 134 2851
rect 94 2802 97 2818
rect 142 2802 145 2848
rect 158 2832 161 2918
rect 238 2872 241 2928
rect 210 2868 214 2871
rect 226 2868 230 2871
rect 270 2862 273 3148
rect 294 3062 297 3148
rect 406 3142 409 3148
rect 422 3122 425 3128
rect 310 3102 313 3118
rect 342 3062 345 3068
rect 310 3031 313 3050
rect 358 3032 361 3078
rect 443 3068 446 3071
rect 454 3052 457 3068
rect 344 3003 346 3007
rect 350 3003 353 3007
rect 357 3003 360 3007
rect 366 2960 369 2979
rect 454 2952 457 3048
rect 310 2932 313 2938
rect 334 2882 337 2938
rect 342 2902 345 2948
rect 218 2858 222 2861
rect 250 2848 254 2851
rect 286 2831 289 2850
rect 318 2832 321 2868
rect 374 2862 377 2868
rect 162 2818 166 2821
rect 182 2762 185 2788
rect 134 2742 137 2748
rect 74 2668 78 2671
rect 62 2492 65 2618
rect 78 2532 81 2668
rect 118 2582 121 2728
rect 174 2662 177 2748
rect 214 2712 217 2718
rect 230 2682 233 2828
rect 294 2732 297 2808
rect 344 2803 346 2807
rect 350 2803 353 2807
rect 357 2803 360 2807
rect 358 2762 361 2788
rect 342 2752 345 2758
rect 310 2742 313 2748
rect 214 2672 217 2678
rect 318 2672 321 2708
rect 374 2692 377 2738
rect 398 2712 401 2938
rect 414 2932 417 2938
rect 414 2812 417 2928
rect 462 2902 465 3538
rect 534 3482 537 3488
rect 550 3412 553 3468
rect 606 3462 609 3548
rect 942 3541 945 3548
rect 934 3538 945 3541
rect 662 3532 665 3538
rect 902 3532 905 3538
rect 646 3492 649 3528
rect 886 3522 889 3528
rect 702 3482 705 3518
rect 848 3503 850 3507
rect 854 3503 857 3507
rect 861 3503 864 3507
rect 886 3501 889 3518
rect 886 3498 897 3501
rect 894 3482 897 3498
rect 602 3458 606 3461
rect 566 3360 569 3379
rect 582 3352 585 3458
rect 630 3452 633 3458
rect 598 3422 601 3448
rect 638 3422 641 3448
rect 518 3322 521 3328
rect 534 3322 537 3338
rect 470 3262 473 3298
rect 478 3272 481 3278
rect 518 3272 521 3288
rect 506 3268 510 3271
rect 534 3252 537 3278
rect 550 3272 553 3308
rect 598 3272 601 3408
rect 646 3392 649 3448
rect 606 3342 609 3358
rect 606 3272 609 3318
rect 614 3272 617 3328
rect 622 3302 625 3338
rect 630 3312 633 3358
rect 646 3302 649 3348
rect 654 3342 657 3398
rect 670 3392 673 3408
rect 654 3272 657 3338
rect 662 3292 665 3318
rect 686 3302 689 3468
rect 742 3352 745 3458
rect 830 3422 833 3448
rect 782 3342 785 3418
rect 830 3360 833 3379
rect 846 3352 849 3458
rect 878 3372 881 3468
rect 934 3462 937 3538
rect 958 3532 961 3628
rect 990 3592 993 3628
rect 1070 3628 1074 3632
rect 1174 3628 1178 3632
rect 1190 3628 1194 3632
rect 1206 3631 1210 3632
rect 1270 3631 1274 3632
rect 1206 3628 1217 3631
rect 1270 3628 1281 3631
rect 1070 3602 1073 3628
rect 1014 3562 1017 3588
rect 782 3322 785 3328
rect 702 3312 705 3318
rect 694 3272 697 3308
rect 554 3268 558 3271
rect 706 3268 710 3271
rect 570 3248 574 3251
rect 478 3062 481 3238
rect 486 3072 489 3208
rect 486 3062 489 3068
rect 478 2872 481 3058
rect 502 3022 505 3118
rect 494 3002 497 3018
rect 510 3011 513 3248
rect 530 3238 534 3241
rect 534 3162 537 3188
rect 582 3182 585 3268
rect 678 3262 681 3268
rect 618 3258 622 3261
rect 602 3248 606 3251
rect 630 3222 633 3258
rect 654 3248 662 3251
rect 530 3148 534 3151
rect 518 3062 521 3148
rect 582 3142 585 3148
rect 518 3052 521 3058
rect 502 3008 513 3011
rect 502 2922 505 3008
rect 526 2992 529 3138
rect 598 3122 601 3128
rect 582 3082 585 3088
rect 566 3072 569 3078
rect 534 3022 537 3050
rect 622 3032 625 3058
rect 654 3031 657 3248
rect 678 3192 681 3198
rect 686 3141 689 3268
rect 694 3202 697 3268
rect 710 3262 713 3268
rect 766 3261 769 3298
rect 774 3272 777 3308
rect 782 3272 785 3278
rect 798 3272 801 3338
rect 830 3272 833 3338
rect 846 3332 849 3348
rect 848 3303 850 3307
rect 854 3303 857 3307
rect 861 3303 864 3307
rect 870 3302 873 3358
rect 886 3352 889 3378
rect 882 3348 886 3351
rect 870 3291 873 3298
rect 866 3288 873 3291
rect 806 3262 809 3268
rect 814 3262 817 3268
rect 766 3258 777 3261
rect 818 3258 825 3261
rect 718 3242 721 3258
rect 758 3252 761 3258
rect 718 3222 721 3228
rect 702 3152 705 3218
rect 750 3172 753 3238
rect 686 3138 694 3141
rect 698 3138 705 3141
rect 714 3138 718 3141
rect 702 3072 705 3138
rect 734 3132 737 3168
rect 766 3162 769 3248
rect 774 3192 777 3258
rect 794 3248 801 3251
rect 798 3192 801 3248
rect 746 3158 750 3161
rect 674 3058 678 3061
rect 682 3048 689 3051
rect 666 3038 670 3041
rect 654 3028 665 3031
rect 590 2988 598 2991
rect 542 2962 545 2968
rect 514 2958 518 2961
rect 550 2952 553 2968
rect 558 2952 561 2958
rect 498 2918 502 2921
rect 526 2912 529 2948
rect 534 2932 537 2938
rect 566 2892 569 2958
rect 574 2952 577 2978
rect 574 2942 577 2948
rect 510 2862 513 2868
rect 458 2858 462 2861
rect 414 2762 417 2788
rect 422 2752 425 2858
rect 366 2682 369 2688
rect 422 2682 425 2718
rect 430 2711 433 2838
rect 478 2831 481 2850
rect 462 2742 465 2778
rect 526 2742 529 2878
rect 478 2732 481 2738
rect 430 2708 441 2711
rect 342 2662 345 2668
rect 398 2662 401 2668
rect 406 2662 409 2668
rect 422 2662 425 2678
rect 430 2672 433 2678
rect 438 2672 441 2708
rect 478 2692 481 2708
rect 518 2692 521 2708
rect 315 2658 318 2661
rect 354 2658 358 2661
rect 386 2658 390 2661
rect 134 2552 137 2618
rect 174 2552 177 2658
rect 182 2631 185 2650
rect 378 2648 382 2651
rect 366 2612 369 2648
rect 344 2603 346 2607
rect 350 2603 353 2607
rect 357 2603 360 2607
rect 390 2592 393 2658
rect 410 2648 414 2651
rect 182 2562 185 2588
rect 358 2562 361 2588
rect 362 2548 366 2551
rect 182 2542 185 2548
rect 254 2542 257 2548
rect 118 2522 121 2528
rect 134 2512 137 2538
rect 294 2532 297 2538
rect 218 2518 222 2521
rect 174 2482 177 2518
rect 30 2472 33 2478
rect 54 2472 57 2478
rect 90 2468 93 2471
rect 26 2458 30 2461
rect 46 2452 49 2458
rect 30 2372 33 2378
rect 22 2282 25 2348
rect 54 2312 57 2458
rect 82 2448 86 2451
rect 62 2442 65 2448
rect 34 2268 38 2271
rect 22 2252 25 2258
rect 6 2242 9 2248
rect 42 2188 46 2191
rect 34 2148 41 2151
rect 6 2142 9 2148
rect 6 2072 9 2078
rect 22 2042 25 2058
rect 30 2052 33 2068
rect 38 2012 41 2148
rect 54 2072 57 2268
rect 62 2062 65 2308
rect 102 2272 105 2478
rect 174 2422 177 2478
rect 190 2462 193 2468
rect 222 2422 225 2450
rect 110 2272 113 2308
rect 110 2262 113 2268
rect 134 2262 137 2268
rect 142 2262 145 2328
rect 158 2322 161 2338
rect 198 2282 201 2418
rect 206 2362 209 2388
rect 238 2352 241 2458
rect 290 2448 294 2451
rect 310 2432 313 2538
rect 410 2528 414 2531
rect 366 2482 369 2488
rect 344 2403 346 2407
rect 350 2403 353 2407
rect 357 2403 360 2407
rect 246 2362 249 2388
rect 210 2348 214 2351
rect 294 2342 297 2368
rect 354 2348 358 2351
rect 310 2312 313 2328
rect 366 2312 369 2478
rect 382 2472 385 2488
rect 438 2472 441 2668
rect 454 2662 457 2668
rect 462 2662 465 2688
rect 542 2672 545 2768
rect 538 2658 542 2661
rect 502 2652 505 2658
rect 510 2652 513 2658
rect 478 2642 481 2648
rect 486 2642 489 2648
rect 498 2638 502 2641
rect 446 2632 449 2638
rect 534 2560 537 2579
rect 446 2462 449 2548
rect 502 2542 505 2548
rect 462 2492 465 2498
rect 434 2458 438 2461
rect 382 2352 385 2458
rect 454 2452 457 2468
rect 414 2422 417 2450
rect 326 2292 329 2308
rect 326 2282 329 2288
rect 198 2272 201 2278
rect 342 2272 345 2278
rect 249 2268 254 2271
rect 206 2262 209 2268
rect 98 2258 102 2261
rect 114 2248 118 2251
rect 130 2248 134 2251
rect 86 2212 89 2218
rect 118 2132 121 2208
rect 182 2162 185 2188
rect 134 2142 137 2148
rect 118 2122 121 2128
rect 82 2068 86 2071
rect 166 2062 169 2148
rect 206 2132 209 2138
rect 206 2082 209 2128
rect 238 2102 241 2258
rect 246 2252 249 2268
rect 382 2262 385 2348
rect 438 2342 441 2438
rect 470 2392 473 2448
rect 446 2382 449 2388
rect 454 2352 457 2358
rect 478 2342 481 2508
rect 486 2482 489 2528
rect 550 2482 553 2808
rect 574 2742 577 2918
rect 590 2792 593 2988
rect 598 2942 601 2948
rect 606 2942 609 2948
rect 602 2878 606 2881
rect 614 2852 617 2948
rect 622 2882 625 3018
rect 662 2992 665 3028
rect 686 2992 689 3048
rect 694 3002 697 3058
rect 710 2992 713 3128
rect 742 3122 745 3148
rect 738 3068 742 3071
rect 746 3058 750 3061
rect 734 3052 737 3058
rect 758 3051 761 3158
rect 774 3152 777 3178
rect 802 3168 806 3171
rect 794 3158 798 3161
rect 766 3092 769 3128
rect 774 3102 777 3128
rect 782 3112 785 3138
rect 774 3072 777 3078
rect 782 3072 785 3108
rect 798 3092 801 3148
rect 822 3142 825 3258
rect 830 3182 833 3258
rect 886 3172 889 3308
rect 882 3168 886 3171
rect 834 3148 838 3151
rect 842 3138 846 3141
rect 822 3092 825 3118
rect 848 3103 850 3107
rect 854 3103 857 3107
rect 861 3103 864 3107
rect 750 3048 761 3051
rect 710 2982 713 2988
rect 638 2972 641 2978
rect 654 2972 657 2978
rect 678 2972 681 2978
rect 630 2962 633 2968
rect 638 2962 641 2968
rect 694 2962 697 2968
rect 646 2922 649 2948
rect 686 2932 689 2948
rect 634 2918 638 2921
rect 630 2892 633 2908
rect 658 2888 662 2891
rect 670 2872 673 2928
rect 694 2892 697 2958
rect 726 2932 729 2948
rect 650 2858 657 2861
rect 563 2738 566 2741
rect 582 2692 585 2718
rect 586 2678 590 2681
rect 566 2662 569 2678
rect 598 2662 601 2848
rect 646 2782 649 2788
rect 610 2768 614 2771
rect 618 2758 622 2761
rect 610 2748 614 2751
rect 622 2742 625 2748
rect 638 2732 641 2738
rect 630 2702 633 2718
rect 630 2672 633 2678
rect 574 2652 577 2658
rect 586 2648 590 2651
rect 574 2642 577 2648
rect 558 2522 561 2638
rect 566 2561 569 2618
rect 614 2592 617 2668
rect 638 2662 641 2668
rect 622 2652 625 2658
rect 646 2622 649 2668
rect 654 2582 657 2858
rect 662 2802 665 2848
rect 662 2762 665 2788
rect 670 2742 673 2868
rect 678 2862 681 2868
rect 690 2858 694 2861
rect 678 2792 681 2838
rect 702 2771 705 2888
rect 718 2862 721 2888
rect 726 2842 729 2848
rect 714 2838 718 2841
rect 718 2772 721 2838
rect 734 2782 737 3048
rect 750 2992 753 3048
rect 766 3042 769 3048
rect 766 3012 769 3038
rect 782 3002 785 3058
rect 798 3052 801 3078
rect 858 3068 862 3071
rect 842 3058 846 3061
rect 806 3052 809 3058
rect 834 3048 838 3051
rect 786 2988 790 2991
rect 746 2968 750 2971
rect 758 2962 761 2978
rect 750 2952 753 2958
rect 770 2948 777 2951
rect 766 2942 769 2948
rect 750 2892 753 2898
rect 774 2882 777 2948
rect 746 2878 750 2881
rect 746 2868 750 2871
rect 766 2862 769 2868
rect 774 2862 777 2868
rect 786 2858 790 2861
rect 798 2852 801 3048
rect 814 2992 817 3048
rect 854 3012 857 3058
rect 810 2968 814 2971
rect 834 2958 841 2961
rect 814 2952 817 2958
rect 830 2952 833 2958
rect 814 2942 817 2948
rect 806 2892 809 2928
rect 742 2792 745 2828
rect 702 2768 713 2771
rect 710 2762 713 2768
rect 694 2758 702 2761
rect 662 2682 665 2728
rect 670 2712 673 2738
rect 678 2701 681 2748
rect 670 2698 681 2701
rect 670 2672 673 2698
rect 694 2692 697 2758
rect 710 2752 713 2758
rect 742 2742 745 2748
rect 730 2738 734 2741
rect 742 2731 745 2738
rect 734 2728 745 2731
rect 710 2702 713 2728
rect 702 2662 705 2668
rect 710 2662 713 2698
rect 726 2662 729 2668
rect 646 2562 649 2568
rect 654 2562 657 2568
rect 566 2558 574 2561
rect 670 2552 673 2578
rect 678 2552 681 2658
rect 722 2648 726 2651
rect 694 2642 697 2648
rect 686 2562 689 2638
rect 734 2632 737 2728
rect 750 2692 753 2848
rect 782 2832 785 2838
rect 798 2822 801 2848
rect 806 2802 809 2848
rect 774 2782 777 2788
rect 806 2782 809 2788
rect 798 2772 801 2778
rect 786 2768 790 2771
rect 758 2762 761 2768
rect 770 2758 774 2761
rect 794 2758 798 2761
rect 806 2752 809 2768
rect 778 2748 782 2751
rect 762 2678 766 2681
rect 746 2668 750 2671
rect 742 2652 745 2658
rect 758 2592 761 2638
rect 766 2622 769 2668
rect 774 2662 777 2688
rect 782 2672 785 2678
rect 798 2672 801 2678
rect 790 2632 793 2658
rect 806 2622 809 2668
rect 814 2662 817 2898
rect 826 2868 830 2871
rect 838 2862 841 2958
rect 850 2948 854 2951
rect 862 2942 865 3008
rect 870 2962 873 3158
rect 878 3152 881 3158
rect 870 2932 873 2938
rect 848 2903 850 2907
rect 854 2903 857 2907
rect 861 2903 864 2907
rect 878 2892 881 2978
rect 894 2972 897 3458
rect 974 3392 977 3548
rect 1014 3462 1017 3548
rect 1062 3532 1065 3538
rect 1078 3532 1081 3568
rect 1154 3548 1159 3551
rect 1118 3542 1121 3548
rect 1078 3512 1081 3528
rect 1166 3512 1169 3548
rect 1174 3501 1177 3628
rect 1190 3592 1193 3628
rect 1214 3592 1217 3628
rect 1278 3592 1281 3628
rect 1334 3628 1338 3632
rect 1382 3628 1386 3632
rect 1422 3631 1426 3632
rect 1446 3631 1450 3632
rect 1422 3628 1433 3631
rect 1446 3628 1457 3631
rect 1334 3602 1337 3628
rect 1360 3603 1362 3607
rect 1366 3603 1369 3607
rect 1373 3603 1376 3607
rect 1238 3562 1241 3588
rect 1382 3582 1385 3628
rect 1430 3592 1433 3628
rect 1454 3592 1457 3628
rect 1462 3628 1466 3632
rect 1478 3628 1482 3632
rect 1510 3628 1514 3632
rect 1526 3628 1530 3632
rect 1574 3628 1578 3632
rect 1606 3628 1610 3632
rect 1662 3628 1666 3632
rect 1694 3628 1698 3632
rect 1718 3631 1722 3632
rect 1718 3628 1729 3631
rect 1462 3602 1465 3628
rect 1478 3592 1481 3628
rect 1510 3602 1513 3628
rect 1526 3592 1529 3628
rect 1574 3602 1577 3628
rect 1606 3602 1609 3628
rect 1506 3588 1510 3591
rect 1542 3560 1545 3579
rect 1202 3548 1206 3551
rect 1387 3548 1390 3551
rect 1466 3548 1470 3551
rect 1238 3542 1241 3548
rect 1166 3498 1177 3501
rect 1166 3492 1169 3498
rect 1230 3492 1233 3518
rect 1286 3512 1289 3538
rect 1302 3522 1305 3528
rect 1302 3492 1305 3508
rect 1342 3492 1345 3548
rect 1350 3492 1353 3538
rect 1398 3512 1401 3548
rect 1438 3502 1441 3548
rect 1486 3542 1489 3548
rect 1274 3488 1278 3491
rect 986 3438 990 3441
rect 1014 3392 1017 3458
rect 1022 3431 1025 3450
rect 1054 3432 1057 3468
rect 902 3322 905 3328
rect 902 3262 905 3318
rect 926 3312 929 3368
rect 946 3358 950 3361
rect 998 3352 1001 3378
rect 1054 3362 1057 3408
rect 1062 3392 1065 3418
rect 938 3348 942 3351
rect 1050 3348 1054 3351
rect 1038 3342 1041 3348
rect 986 3338 990 3341
rect 1026 3338 1030 3341
rect 942 3272 945 3278
rect 958 3272 961 3338
rect 974 3332 977 3338
rect 982 3302 985 3328
rect 1070 3322 1073 3478
rect 1218 3468 1222 3471
rect 1238 3462 1241 3478
rect 1274 3468 1278 3471
rect 1306 3468 1310 3471
rect 1210 3458 1214 3461
rect 1090 3388 1094 3391
rect 1110 3352 1113 3458
rect 1222 3452 1225 3458
rect 1190 3432 1193 3448
rect 1154 3428 1158 3431
rect 1246 3402 1249 3468
rect 1374 3462 1377 3488
rect 1438 3482 1441 3488
rect 1422 3462 1425 3468
rect 1478 3462 1481 3468
rect 1526 3462 1529 3548
rect 1574 3532 1577 3538
rect 1590 3532 1593 3568
rect 1662 3552 1665 3628
rect 1694 3591 1697 3628
rect 1726 3592 1729 3628
rect 1758 3628 1762 3632
rect 1774 3631 1778 3632
rect 1766 3628 1778 3631
rect 1790 3628 1794 3632
rect 1902 3628 1906 3632
rect 1934 3631 1938 3632
rect 1958 3631 1962 3632
rect 1934 3628 1945 3631
rect 1758 3602 1761 3628
rect 1694 3588 1702 3591
rect 1750 3562 1753 3588
rect 1630 3532 1633 3548
rect 1710 3482 1713 3548
rect 1750 3532 1753 3548
rect 1766 3531 1769 3628
rect 1790 3592 1793 3628
rect 1902 3602 1905 3628
rect 1942 3592 1945 3628
rect 1950 3628 1962 3631
rect 1974 3628 1978 3632
rect 2062 3628 2066 3632
rect 2078 3628 2082 3632
rect 2118 3628 2122 3632
rect 2230 3628 2234 3632
rect 2406 3628 2410 3632
rect 1950 3592 1953 3628
rect 1974 3602 1977 3628
rect 2062 3572 2065 3628
rect 2078 3592 2081 3628
rect 2230 3602 2233 3628
rect 2384 3603 2386 3607
rect 2390 3603 2393 3607
rect 2397 3603 2400 3607
rect 2406 3602 2409 3628
rect 3408 3603 3410 3607
rect 3414 3603 3417 3607
rect 3421 3603 3424 3607
rect 2230 3560 2233 3579
rect 1758 3528 1769 3531
rect 1798 3532 1801 3538
rect 1814 3532 1817 3538
rect 1614 3472 1617 3478
rect 1258 3458 1262 3461
rect 1314 3458 1318 3461
rect 1546 3458 1550 3461
rect 1262 3448 1270 3451
rect 1262 3442 1265 3448
rect 1130 3348 1134 3351
rect 1086 3302 1089 3348
rect 1190 3332 1193 3338
rect 1110 3272 1113 3278
rect 1094 3262 1097 3268
rect 1042 3258 1046 3261
rect 1014 3252 1017 3258
rect 990 3231 993 3250
rect 1062 3231 1065 3250
rect 922 3168 926 3171
rect 966 3152 969 3208
rect 1166 3192 1169 3218
rect 1174 3192 1177 3328
rect 1190 3292 1193 3318
rect 1230 3292 1233 3368
rect 1238 3362 1241 3388
rect 1262 3352 1265 3438
rect 1270 3392 1273 3418
rect 1238 3292 1241 3348
rect 1270 3342 1273 3348
rect 1238 3282 1241 3288
rect 1262 3282 1265 3338
rect 1286 3312 1289 3458
rect 1302 3392 1305 3448
rect 1310 3362 1313 3368
rect 1294 3352 1297 3358
rect 1306 3348 1310 3351
rect 1318 3331 1321 3428
rect 1326 3342 1329 3348
rect 1318 3328 1326 3331
rect 1326 3302 1329 3328
rect 1334 3292 1337 3448
rect 1390 3431 1393 3450
rect 1518 3432 1521 3438
rect 1360 3403 1362 3407
rect 1366 3403 1369 3407
rect 1373 3403 1376 3407
rect 1206 3272 1209 3278
rect 1342 3272 1345 3398
rect 1402 3388 1406 3391
rect 1370 3358 1374 3361
rect 1362 3348 1366 3351
rect 1350 3342 1353 3348
rect 1198 3268 1206 3271
rect 1306 3268 1310 3271
rect 1322 3268 1326 3271
rect 982 3162 985 3168
rect 1002 3158 1006 3161
rect 1038 3160 1041 3179
rect 970 3148 974 3151
rect 1018 3148 1022 3151
rect 918 3142 921 3148
rect 906 3138 910 3141
rect 938 3138 942 3141
rect 958 3141 961 3148
rect 982 3142 985 3148
rect 958 3138 974 3141
rect 938 3128 942 3131
rect 910 3082 913 3118
rect 966 3082 969 3088
rect 950 3062 953 3068
rect 1006 3062 1009 3148
rect 1126 3142 1129 3148
rect 1050 3078 1054 3081
rect 1070 3072 1073 3138
rect 1086 3102 1089 3128
rect 1094 3108 1102 3111
rect 1094 3092 1097 3108
rect 1134 3072 1137 3078
rect 1082 3068 1086 3071
rect 1114 3068 1118 3071
rect 1134 3062 1137 3068
rect 902 3032 905 3058
rect 918 3031 921 3050
rect 918 2992 921 2998
rect 914 2968 918 2971
rect 858 2868 862 2871
rect 886 2862 889 2918
rect 822 2752 825 2858
rect 854 2852 857 2858
rect 838 2842 841 2848
rect 854 2812 857 2818
rect 838 2762 841 2768
rect 862 2762 865 2858
rect 878 2762 881 2818
rect 838 2742 841 2748
rect 886 2742 889 2848
rect 894 2812 897 2968
rect 938 2958 942 2961
rect 918 2952 921 2958
rect 902 2862 905 2928
rect 934 2922 937 2938
rect 910 2872 913 2918
rect 934 2892 937 2918
rect 950 2912 953 2948
rect 958 2942 961 2998
rect 1006 2992 1009 3048
rect 1062 3042 1065 3048
rect 1078 3042 1081 3058
rect 1110 3052 1113 3058
rect 1090 3048 1094 3051
rect 966 2972 969 2978
rect 1002 2968 1006 2971
rect 978 2958 982 2961
rect 978 2938 982 2941
rect 974 2928 982 2931
rect 910 2862 913 2868
rect 918 2862 921 2878
rect 902 2762 905 2858
rect 918 2792 921 2858
rect 950 2852 953 2908
rect 974 2862 977 2928
rect 1006 2922 1009 2948
rect 986 2888 990 2891
rect 998 2872 1001 2888
rect 1014 2872 1017 2958
rect 1030 2872 1033 3028
rect 1078 3002 1081 3038
rect 1110 3032 1113 3048
rect 1134 3042 1137 3048
rect 1126 3012 1129 3018
rect 1038 2962 1041 2988
rect 1142 2952 1145 3148
rect 1190 3142 1193 3218
rect 1198 3132 1201 3268
rect 1262 3262 1265 3268
rect 1286 3262 1289 3268
rect 1218 3258 1222 3261
rect 1234 3258 1238 3261
rect 1298 3258 1302 3261
rect 1258 3248 1262 3251
rect 1230 3232 1233 3248
rect 1262 3232 1265 3238
rect 1270 3232 1273 3238
rect 1302 3202 1305 3258
rect 1214 3162 1217 3188
rect 1210 3148 1214 3151
rect 1158 3118 1166 3121
rect 1158 3072 1161 3118
rect 1182 3052 1185 3118
rect 1170 3028 1174 3031
rect 1086 2932 1089 2938
rect 962 2818 966 2821
rect 926 2772 929 2778
rect 942 2762 945 2768
rect 830 2732 833 2738
rect 830 2692 833 2708
rect 848 2703 850 2707
rect 854 2703 857 2707
rect 861 2703 864 2707
rect 878 2702 881 2718
rect 894 2692 897 2748
rect 910 2742 913 2758
rect 926 2752 929 2758
rect 902 2722 905 2738
rect 926 2702 929 2748
rect 942 2742 945 2748
rect 974 2742 977 2858
rect 982 2792 985 2848
rect 1006 2842 1009 2848
rect 1022 2812 1025 2858
rect 1030 2762 1033 2868
rect 1054 2862 1057 2918
rect 1094 2872 1097 2878
rect 1074 2858 1078 2861
rect 1046 2832 1049 2838
rect 1046 2792 1049 2808
rect 990 2758 998 2761
rect 990 2752 993 2758
rect 1014 2752 1017 2758
rect 954 2738 958 2741
rect 934 2732 937 2738
rect 990 2732 993 2738
rect 958 2728 966 2731
rect 850 2688 854 2691
rect 862 2672 865 2678
rect 918 2672 921 2688
rect 926 2682 929 2698
rect 950 2692 953 2728
rect 958 2712 961 2728
rect 998 2722 1001 2748
rect 1030 2742 1033 2748
rect 1022 2732 1025 2738
rect 1046 2722 1049 2728
rect 966 2692 969 2708
rect 974 2682 977 2688
rect 954 2668 958 2671
rect 830 2632 833 2658
rect 838 2592 841 2668
rect 918 2662 921 2668
rect 946 2658 950 2661
rect 902 2652 905 2658
rect 846 2612 849 2638
rect 894 2632 897 2638
rect 826 2588 830 2591
rect 694 2562 697 2578
rect 706 2568 710 2571
rect 762 2568 766 2571
rect 722 2558 726 2561
rect 574 2542 577 2548
rect 630 2542 633 2548
rect 670 2538 678 2541
rect 598 2482 601 2538
rect 606 2532 609 2538
rect 622 2512 625 2538
rect 630 2502 633 2538
rect 638 2492 641 2538
rect 534 2462 537 2468
rect 494 2452 497 2458
rect 486 2422 489 2448
rect 494 2392 497 2428
rect 550 2402 553 2478
rect 635 2468 638 2471
rect 654 2462 657 2518
rect 670 2492 673 2538
rect 686 2512 689 2558
rect 738 2548 742 2551
rect 702 2541 705 2548
rect 702 2538 718 2541
rect 738 2538 742 2541
rect 710 2492 713 2518
rect 750 2512 753 2558
rect 758 2552 761 2558
rect 782 2542 785 2588
rect 826 2568 830 2571
rect 794 2558 798 2561
rect 794 2548 798 2551
rect 782 2532 785 2538
rect 806 2522 809 2558
rect 814 2512 817 2558
rect 826 2548 830 2551
rect 846 2542 849 2608
rect 862 2542 865 2598
rect 870 2552 873 2598
rect 886 2572 889 2618
rect 902 2592 905 2608
rect 890 2558 894 2561
rect 882 2548 886 2551
rect 866 2538 873 2541
rect 646 2442 649 2448
rect 558 2382 561 2388
rect 486 2352 489 2378
rect 526 2372 529 2378
rect 542 2362 545 2368
rect 590 2362 593 2408
rect 598 2362 601 2438
rect 606 2372 609 2378
rect 614 2372 617 2378
rect 514 2358 518 2361
rect 610 2348 614 2351
rect 482 2338 486 2341
rect 430 2332 433 2338
rect 390 2262 393 2318
rect 446 2272 449 2338
rect 486 2292 489 2298
rect 462 2272 465 2278
rect 418 2268 422 2271
rect 390 2222 393 2248
rect 344 2203 346 2207
rect 350 2203 353 2207
rect 357 2203 360 2207
rect 326 2160 329 2179
rect 358 2142 361 2158
rect 418 2148 422 2151
rect 374 2122 377 2128
rect 262 2082 265 2118
rect 398 2092 401 2108
rect 438 2102 441 2218
rect 398 2082 401 2088
rect 446 2082 449 2268
rect 470 2212 473 2248
rect 478 2192 481 2258
rect 494 2152 497 2348
rect 514 2338 518 2341
rect 526 2332 529 2348
rect 562 2338 566 2341
rect 550 2302 553 2338
rect 522 2258 526 2261
rect 566 2182 569 2278
rect 582 2272 585 2338
rect 614 2231 617 2250
rect 590 2192 593 2208
rect 622 2192 625 2358
rect 630 2192 633 2418
rect 638 2392 641 2438
rect 654 2412 657 2418
rect 670 2392 673 2488
rect 710 2471 713 2478
rect 710 2468 718 2471
rect 678 2462 681 2468
rect 686 2462 689 2468
rect 638 2382 641 2388
rect 682 2368 686 2371
rect 670 2362 673 2368
rect 694 2352 697 2458
rect 702 2362 705 2448
rect 658 2348 662 2351
rect 662 2292 665 2338
rect 678 2332 681 2338
rect 686 2332 689 2348
rect 710 2342 713 2468
rect 730 2458 734 2461
rect 746 2458 750 2461
rect 770 2458 774 2461
rect 782 2452 785 2508
rect 798 2478 806 2481
rect 790 2452 793 2458
rect 782 2442 785 2448
rect 766 2381 769 2438
rect 762 2378 769 2381
rect 790 2422 793 2438
rect 758 2372 761 2378
rect 718 2352 721 2358
rect 742 2352 745 2358
rect 754 2348 758 2351
rect 718 2342 721 2348
rect 774 2342 777 2368
rect 790 2362 793 2418
rect 798 2352 801 2478
rect 806 2472 809 2478
rect 810 2458 814 2461
rect 822 2451 825 2518
rect 870 2512 873 2538
rect 886 2538 894 2541
rect 848 2503 850 2507
rect 854 2503 857 2507
rect 861 2503 864 2507
rect 834 2468 838 2471
rect 886 2462 889 2538
rect 894 2462 897 2468
rect 818 2448 825 2451
rect 834 2458 838 2461
rect 830 2372 833 2458
rect 870 2442 873 2448
rect 838 2392 841 2428
rect 826 2358 830 2361
rect 818 2348 822 2351
rect 862 2342 865 2368
rect 886 2352 889 2458
rect 902 2451 905 2458
rect 894 2448 905 2451
rect 910 2452 913 2648
rect 918 2612 921 2658
rect 918 2542 921 2548
rect 918 2462 921 2528
rect 926 2492 929 2658
rect 958 2651 961 2658
rect 946 2648 961 2651
rect 982 2632 985 2668
rect 990 2662 993 2678
rect 998 2672 1001 2688
rect 1030 2682 1033 2688
rect 1046 2682 1049 2708
rect 1054 2692 1057 2848
rect 1086 2842 1089 2858
rect 1062 2742 1065 2748
rect 1006 2632 1009 2658
rect 1014 2632 1017 2668
rect 1038 2662 1041 2668
rect 1026 2658 1030 2661
rect 974 2592 977 2598
rect 1046 2592 1049 2598
rect 934 2582 937 2588
rect 954 2548 958 2551
rect 974 2492 977 2568
rect 1006 2562 1009 2568
rect 986 2548 990 2551
rect 1006 2502 1009 2558
rect 1054 2552 1057 2648
rect 1062 2612 1065 2718
rect 1070 2662 1073 2818
rect 1094 2742 1097 2748
rect 1078 2702 1081 2718
rect 1082 2678 1086 2681
rect 1082 2668 1086 2671
rect 1062 2542 1065 2608
rect 1078 2602 1081 2668
rect 1086 2592 1089 2628
rect 1078 2552 1081 2558
rect 1094 2552 1097 2738
rect 1102 2672 1105 2928
rect 1142 2912 1145 2948
rect 1198 2942 1201 3128
rect 1206 3062 1209 3148
rect 1262 3142 1265 3148
rect 1278 3132 1281 3188
rect 1318 3142 1321 3268
rect 1350 3262 1353 3308
rect 1374 3292 1377 3348
rect 1334 3252 1337 3258
rect 1362 3248 1366 3251
rect 1246 3082 1249 3098
rect 1334 3092 1337 3228
rect 1360 3203 1362 3207
rect 1366 3203 1369 3207
rect 1373 3203 1376 3207
rect 1262 3072 1265 3078
rect 1294 3031 1297 3050
rect 1330 3048 1334 3051
rect 1262 2972 1265 2978
rect 1222 2962 1225 2968
rect 1230 2962 1233 2968
rect 1278 2962 1281 2988
rect 1294 2972 1297 2978
rect 1318 2972 1321 2978
rect 1206 2952 1209 2958
rect 1286 2952 1289 2968
rect 1306 2958 1310 2961
rect 1318 2952 1321 2958
rect 1246 2942 1249 2948
rect 1342 2942 1345 3198
rect 1382 3172 1385 3288
rect 1350 3072 1353 3088
rect 1382 3072 1385 3168
rect 1378 3058 1382 3061
rect 1390 3052 1393 3318
rect 1398 3292 1401 3318
rect 1422 3292 1425 3338
rect 1478 3332 1481 3378
rect 1526 3352 1529 3458
rect 1566 3422 1569 3450
rect 1582 3392 1585 3398
rect 1542 3362 1545 3388
rect 1598 3372 1601 3468
rect 1606 3418 1614 3421
rect 1606 3372 1609 3418
rect 1718 3402 1721 3418
rect 1742 3392 1745 3478
rect 1622 3382 1625 3388
rect 1742 3382 1745 3388
rect 1590 3362 1593 3368
rect 1562 3348 1566 3351
rect 1594 3338 1598 3341
rect 1494 3332 1497 3338
rect 1590 3322 1593 3338
rect 1462 3282 1465 3288
rect 1406 3262 1409 3278
rect 1446 3252 1449 3268
rect 1478 3262 1481 3318
rect 1510 3292 1513 3308
rect 1486 3272 1489 3278
rect 1490 3248 1494 3251
rect 1398 3242 1401 3248
rect 1398 3212 1401 3238
rect 1406 3142 1409 3248
rect 1414 3162 1417 3248
rect 1454 3172 1457 3208
rect 1494 3162 1497 3168
rect 1502 3162 1505 3288
rect 1606 3272 1609 3328
rect 1510 3192 1513 3248
rect 1526 3232 1529 3258
rect 1542 3242 1545 3248
rect 1518 3162 1521 3168
rect 1526 3162 1529 3178
rect 1538 3168 1542 3171
rect 1434 3158 1438 3161
rect 1426 3148 1430 3151
rect 1450 3148 1454 3151
rect 1490 3148 1494 3151
rect 1414 3142 1417 3148
rect 1466 3138 1470 3141
rect 1406 3132 1409 3138
rect 1478 3132 1481 3148
rect 1438 3072 1441 3128
rect 1454 3072 1457 3078
rect 1470 3062 1473 3078
rect 1478 3072 1481 3078
rect 1450 3058 1454 3061
rect 1466 3058 1470 3061
rect 1402 3048 1406 3051
rect 1218 2938 1222 2941
rect 1306 2938 1310 2941
rect 1230 2932 1233 2938
rect 1186 2928 1190 2931
rect 1350 2931 1353 3048
rect 1360 3003 1362 3007
rect 1366 3003 1369 3007
rect 1373 3003 1376 3007
rect 1370 2968 1374 2971
rect 1382 2962 1385 3018
rect 1342 2928 1353 2931
rect 1110 2792 1113 2908
rect 1126 2862 1129 2908
rect 1182 2872 1185 2878
rect 1310 2872 1313 2878
rect 1267 2868 1270 2871
rect 1290 2868 1294 2871
rect 1166 2862 1169 2868
rect 1134 2822 1137 2850
rect 1130 2788 1134 2791
rect 1222 2791 1225 2858
rect 1270 2842 1273 2848
rect 1294 2822 1297 2848
rect 1222 2788 1233 2791
rect 1110 2782 1113 2788
rect 1110 2692 1113 2758
rect 1230 2752 1233 2788
rect 1278 2762 1281 2788
rect 1214 2732 1217 2738
rect 1230 2732 1233 2738
rect 1294 2722 1297 2818
rect 1302 2802 1305 2818
rect 1318 2742 1321 2808
rect 1326 2752 1329 2908
rect 1334 2892 1337 2898
rect 1334 2862 1337 2888
rect 1342 2852 1345 2928
rect 1366 2902 1369 2918
rect 1350 2882 1353 2898
rect 1354 2868 1358 2871
rect 1366 2852 1369 2868
rect 1338 2848 1342 2851
rect 1334 2832 1337 2838
rect 1342 2832 1345 2838
rect 1334 2762 1337 2768
rect 1342 2752 1345 2828
rect 1382 2812 1385 2858
rect 1390 2832 1393 3038
rect 1414 3022 1417 3058
rect 1430 3052 1433 3058
rect 1462 3042 1465 3048
rect 1422 3032 1425 3038
rect 1446 2992 1449 3028
rect 1486 2992 1489 3068
rect 1502 3062 1505 3158
rect 1526 3142 1529 3158
rect 1550 3142 1553 3238
rect 1514 3138 1518 3141
rect 1542 3138 1550 3141
rect 1542 3112 1545 3138
rect 1522 3088 1526 3091
rect 1530 3068 1534 3071
rect 1550 3062 1553 3088
rect 1558 3062 1561 3208
rect 1606 3192 1609 3268
rect 1614 3182 1617 3218
rect 1614 3162 1617 3178
rect 1574 3072 1577 3078
rect 1582 3062 1585 3138
rect 1610 3118 1614 3121
rect 1622 3092 1625 3368
rect 1750 3352 1753 3528
rect 1758 3352 1761 3528
rect 1798 3392 1801 3478
rect 1814 3472 1817 3478
rect 1846 3422 1849 3450
rect 1854 3422 1857 3528
rect 1880 3503 1882 3507
rect 1886 3503 1889 3507
rect 1893 3503 1896 3507
rect 1902 3472 1905 3508
rect 1966 3502 1969 3548
rect 1990 3542 1993 3548
rect 1998 3542 2001 3548
rect 2022 3542 2025 3558
rect 2162 3538 2166 3541
rect 2014 3532 2017 3538
rect 1974 3522 1977 3528
rect 1982 3512 1985 3518
rect 2038 3502 2041 3518
rect 1862 3442 1865 3458
rect 1910 3402 1913 3418
rect 1950 3392 1953 3498
rect 2038 3492 2041 3498
rect 2094 3492 2097 3538
rect 2190 3532 2193 3548
rect 2170 3528 2174 3531
rect 2174 3522 2177 3528
rect 2182 3492 2185 3518
rect 1990 3482 1993 3488
rect 2006 3462 2009 3468
rect 2046 3442 2049 3458
rect 2046 3411 2049 3438
rect 2054 3422 2057 3448
rect 2046 3408 2057 3411
rect 1822 3360 1825 3379
rect 1986 3358 1990 3361
rect 1802 3348 1806 3351
rect 1678 3332 1681 3338
rect 1758 3302 1761 3348
rect 1778 3338 1782 3341
rect 1782 3322 1785 3338
rect 1854 3332 1857 3338
rect 1694 3282 1697 3298
rect 1870 3292 1873 3328
rect 1974 3322 1977 3358
rect 1998 3342 2001 3358
rect 1880 3303 1882 3307
rect 1886 3303 1889 3307
rect 1893 3303 1896 3307
rect 1630 3262 1633 3278
rect 1638 3262 1641 3268
rect 1662 3262 1665 3278
rect 1674 3268 1678 3271
rect 1646 3161 1649 3218
rect 1686 3162 1689 3278
rect 1694 3262 1697 3278
rect 1646 3158 1657 3161
rect 1654 3152 1657 3158
rect 1686 3152 1689 3158
rect 1642 3148 1646 3151
rect 1630 3122 1633 3128
rect 1598 3082 1601 3088
rect 1614 3062 1617 3088
rect 1630 3082 1633 3118
rect 1538 3058 1542 3061
rect 1498 3048 1502 3051
rect 1406 2942 1409 2948
rect 1438 2942 1441 2948
rect 1446 2942 1449 2978
rect 1474 2958 1478 2961
rect 1398 2922 1401 2938
rect 1422 2932 1425 2938
rect 1410 2878 1422 2881
rect 1434 2868 1438 2871
rect 1398 2842 1401 2848
rect 1360 2803 1362 2807
rect 1366 2803 1369 2807
rect 1373 2803 1376 2807
rect 1406 2762 1409 2828
rect 1414 2792 1417 2868
rect 1422 2862 1425 2868
rect 1446 2862 1449 2868
rect 1454 2852 1457 2958
rect 1486 2952 1489 2968
rect 1462 2932 1465 2938
rect 1462 2892 1465 2918
rect 1470 2872 1473 2948
rect 1494 2941 1497 2968
rect 1526 2962 1529 3058
rect 1542 2992 1545 3048
rect 1558 3042 1561 3058
rect 1550 3032 1553 3038
rect 1574 2992 1577 2998
rect 1582 2992 1585 3058
rect 1638 3052 1641 3058
rect 1594 3048 1598 3051
rect 1606 3032 1609 3048
rect 1626 3038 1630 3041
rect 1578 2968 1582 2971
rect 1558 2962 1561 2968
rect 1622 2962 1625 2968
rect 1610 2958 1614 2961
rect 1486 2938 1497 2941
rect 1514 2938 1518 2941
rect 1470 2852 1473 2858
rect 1454 2832 1457 2848
rect 1486 2842 1489 2938
rect 1534 2922 1537 2948
rect 1546 2938 1550 2941
rect 1494 2872 1497 2878
rect 1510 2872 1513 2878
rect 1454 2792 1457 2798
rect 1470 2772 1473 2838
rect 1526 2832 1529 2918
rect 1486 2792 1489 2818
rect 1418 2768 1422 2771
rect 1366 2752 1369 2758
rect 1398 2742 1401 2748
rect 1406 2742 1409 2758
rect 1466 2748 1470 2751
rect 1102 2632 1105 2658
rect 1118 2582 1121 2718
rect 1146 2688 1150 2691
rect 1126 2672 1129 2678
rect 1118 2562 1121 2578
rect 1134 2542 1137 2548
rect 1098 2538 1102 2541
rect 946 2488 950 2491
rect 1006 2488 1014 2491
rect 934 2472 937 2488
rect 998 2482 1001 2488
rect 962 2468 966 2471
rect 994 2468 998 2471
rect 894 2352 897 2448
rect 914 2428 918 2431
rect 910 2352 913 2388
rect 926 2362 929 2468
rect 938 2458 942 2461
rect 954 2458 958 2461
rect 706 2338 710 2341
rect 802 2338 806 2341
rect 882 2338 886 2341
rect 790 2332 793 2338
rect 678 2272 681 2328
rect 734 2302 737 2318
rect 742 2282 745 2308
rect 758 2272 761 2298
rect 838 2262 841 2318
rect 894 2312 897 2348
rect 918 2342 921 2358
rect 926 2342 929 2348
rect 902 2322 905 2338
rect 934 2332 937 2338
rect 848 2303 850 2307
rect 854 2303 857 2307
rect 861 2303 864 2307
rect 926 2292 929 2308
rect 698 2258 702 2261
rect 858 2258 862 2261
rect 898 2258 902 2261
rect 638 2252 641 2258
rect 598 2172 601 2178
rect 630 2172 633 2178
rect 554 2168 558 2171
rect 526 2162 529 2168
rect 462 2142 465 2148
rect 454 2132 457 2138
rect 222 2072 225 2078
rect 414 2072 417 2078
rect 270 2062 273 2068
rect 358 2062 361 2068
rect 462 2062 465 2138
rect 90 2058 94 2061
rect 321 2058 326 2061
rect 54 2051 57 2058
rect 54 2048 62 2051
rect 82 2048 86 2051
rect 94 2032 97 2038
rect 130 2018 134 2021
rect 10 1988 14 1991
rect 30 1972 33 1978
rect 66 1958 70 1961
rect 22 1952 25 1958
rect 222 1952 225 2058
rect 318 2052 321 2058
rect 254 2022 257 2050
rect 446 2031 449 2050
rect 270 1992 273 2008
rect 238 1962 241 1988
rect 286 1962 289 1968
rect 42 1948 46 1951
rect 66 1948 70 1951
rect 258 1948 262 1951
rect 54 1942 57 1948
rect 294 1942 297 2018
rect 344 2003 346 2007
rect 350 2003 353 2007
rect 357 2003 360 2007
rect 310 1942 313 1948
rect 266 1938 270 1941
rect 190 1932 193 1938
rect 318 1932 321 1998
rect 378 1968 382 1971
rect 174 1922 177 1928
rect 30 1892 33 1908
rect 94 1902 97 1918
rect 134 1872 137 1878
rect 150 1872 153 1878
rect 222 1872 225 1898
rect 202 1858 206 1861
rect 182 1822 185 1850
rect 182 1762 185 1788
rect 206 1752 209 1858
rect 246 1852 249 1858
rect 230 1792 233 1818
rect 186 1748 190 1751
rect 6 1742 9 1748
rect 134 1732 137 1738
rect 118 1722 121 1728
rect 94 1672 97 1678
rect 110 1662 113 1668
rect 206 1662 209 1748
rect 214 1672 217 1718
rect 262 1682 265 1918
rect 302 1902 305 1918
rect 318 1882 321 1928
rect 334 1912 337 1948
rect 358 1942 361 1968
rect 366 1882 369 1918
rect 302 1852 305 1868
rect 362 1858 366 1861
rect 270 1831 273 1850
rect 344 1803 346 1807
rect 350 1803 353 1807
rect 357 1803 360 1807
rect 322 1768 326 1771
rect 326 1752 329 1758
rect 358 1752 361 1758
rect 298 1748 302 1751
rect 338 1748 342 1751
rect 310 1742 313 1748
rect 270 1712 273 1738
rect 334 1732 337 1738
rect 282 1728 286 1731
rect 354 1728 358 1731
rect 366 1682 369 1768
rect 246 1672 249 1678
rect 162 1658 166 1661
rect 142 1622 145 1650
rect 18 1618 25 1621
rect 10 1588 14 1591
rect 22 1552 25 1618
rect 30 1572 33 1578
rect 142 1562 145 1588
rect 158 1552 161 1658
rect 214 1622 217 1650
rect 46 1502 49 1548
rect 190 1542 193 1578
rect 122 1538 126 1541
rect 62 1512 65 1518
rect 86 1482 89 1508
rect 158 1492 161 1538
rect 206 1492 209 1528
rect 262 1512 265 1678
rect 302 1662 305 1668
rect 366 1662 369 1668
rect 298 1558 302 1561
rect 322 1558 326 1561
rect 322 1538 326 1541
rect 290 1528 294 1531
rect 14 1292 17 1448
rect 70 1412 73 1468
rect 126 1431 129 1458
rect 46 1382 49 1388
rect 34 1338 38 1341
rect 158 1332 161 1488
rect 262 1482 265 1488
rect 302 1472 305 1498
rect 206 1452 209 1458
rect 246 1452 249 1468
rect 198 1422 201 1448
rect 170 1418 174 1421
rect 174 1332 177 1338
rect 30 1262 33 1318
rect 118 1292 121 1318
rect 38 1272 41 1278
rect 158 1272 161 1328
rect 106 1268 110 1271
rect 170 1268 174 1271
rect 34 1258 41 1261
rect 6 1042 9 1048
rect 14 992 17 1158
rect 30 1072 33 1078
rect 26 1058 30 1061
rect 38 1051 41 1258
rect 182 1242 185 1278
rect 206 1272 209 1448
rect 254 1392 257 1408
rect 222 1362 225 1388
rect 270 1362 273 1368
rect 278 1352 281 1358
rect 238 1348 246 1351
rect 222 1332 225 1348
rect 238 1331 241 1348
rect 254 1341 257 1348
rect 250 1338 257 1341
rect 294 1342 297 1368
rect 238 1328 249 1331
rect 246 1292 249 1328
rect 222 1252 225 1258
rect 118 1202 121 1218
rect 70 1152 73 1178
rect 70 1132 73 1138
rect 86 1132 89 1198
rect 206 1172 209 1238
rect 214 1192 217 1248
rect 230 1241 233 1258
rect 222 1238 233 1241
rect 254 1252 257 1338
rect 270 1272 273 1288
rect 222 1192 225 1238
rect 254 1222 257 1248
rect 250 1188 254 1191
rect 262 1162 265 1218
rect 278 1172 281 1318
rect 302 1292 305 1468
rect 310 1362 313 1518
rect 178 1148 182 1151
rect 290 1148 294 1151
rect 134 1082 137 1088
rect 190 1082 193 1118
rect 222 1112 225 1148
rect 254 1132 257 1138
rect 238 1092 241 1128
rect 246 1081 249 1118
rect 262 1112 265 1148
rect 278 1132 281 1148
rect 302 1142 305 1248
rect 326 1162 329 1518
rect 334 1382 337 1658
rect 346 1628 350 1631
rect 344 1603 346 1607
rect 350 1603 353 1607
rect 357 1603 360 1607
rect 342 1542 345 1548
rect 366 1542 369 1658
rect 374 1481 377 1868
rect 382 1581 385 1718
rect 390 1682 393 1968
rect 478 1952 481 2118
rect 486 2062 489 2068
rect 494 2042 497 2148
rect 518 2142 521 2148
rect 502 2132 505 2138
rect 502 2092 505 2128
rect 510 2122 513 2128
rect 502 2072 505 2078
rect 522 2068 526 2071
rect 542 2062 545 2158
rect 510 1992 513 2058
rect 526 2012 529 2048
rect 526 1962 529 1988
rect 462 1922 465 1928
rect 406 1862 409 1868
rect 402 1818 406 1821
rect 438 1772 441 1778
rect 446 1762 449 1908
rect 462 1872 465 1908
rect 470 1862 473 1878
rect 478 1872 481 1938
rect 494 1872 497 1898
rect 518 1892 521 1958
rect 534 1872 537 2048
rect 550 2042 553 2168
rect 586 2158 590 2161
rect 618 2158 622 2161
rect 566 2152 569 2158
rect 574 2151 577 2158
rect 574 2148 585 2151
rect 566 2072 569 2118
rect 582 2072 585 2148
rect 626 2148 630 2151
rect 590 2132 593 2148
rect 638 2092 641 2238
rect 662 2222 665 2228
rect 646 2092 649 2128
rect 654 2082 657 2118
rect 542 1961 545 2018
rect 574 2002 577 2058
rect 598 2052 601 2078
rect 626 2058 630 2061
rect 590 2042 593 2048
rect 598 2032 601 2048
rect 542 1958 550 1961
rect 554 1948 558 1951
rect 566 1942 569 1948
rect 574 1942 577 1978
rect 582 1942 585 2018
rect 590 1992 593 2028
rect 550 1881 553 1938
rect 582 1912 585 1938
rect 590 1902 593 1948
rect 550 1878 558 1881
rect 550 1872 553 1878
rect 566 1862 569 1878
rect 590 1872 593 1888
rect 598 1862 601 1998
rect 646 1981 649 2048
rect 654 1992 657 2008
rect 646 1978 657 1981
rect 634 1968 638 1971
rect 642 1958 646 1961
rect 606 1872 609 1878
rect 458 1858 462 1861
rect 546 1858 550 1861
rect 614 1861 617 1958
rect 626 1948 630 1951
rect 622 1872 625 1918
rect 646 1892 649 1948
rect 654 1941 657 1978
rect 662 1972 665 2178
rect 682 2148 686 2151
rect 670 2072 673 2098
rect 670 2012 673 2058
rect 678 1962 681 2038
rect 694 2022 697 2118
rect 702 2062 705 2258
rect 910 2252 913 2258
rect 790 2231 793 2250
rect 758 2192 761 2208
rect 714 2168 718 2171
rect 778 2168 782 2171
rect 738 2158 742 2161
rect 802 2158 806 2161
rect 758 2152 761 2158
rect 822 2152 825 2188
rect 838 2182 841 2218
rect 862 2192 865 2198
rect 886 2152 889 2218
rect 722 2148 726 2151
rect 794 2148 798 2151
rect 762 2138 766 2141
rect 826 2138 830 2141
rect 758 2082 761 2108
rect 806 2072 809 2118
rect 814 2112 817 2128
rect 742 2062 745 2068
rect 798 2052 801 2058
rect 710 2022 713 2050
rect 734 2018 742 2021
rect 694 1972 697 2008
rect 710 1992 713 2008
rect 682 1958 686 1961
rect 694 1952 697 1968
rect 666 1948 670 1951
rect 674 1948 678 1951
rect 694 1942 697 1948
rect 702 1942 705 1988
rect 722 1948 726 1951
rect 654 1938 665 1941
rect 662 1892 665 1938
rect 678 1882 681 1938
rect 722 1928 726 1931
rect 702 1892 705 1928
rect 678 1872 681 1878
rect 710 1872 713 1918
rect 734 1892 737 2018
rect 798 2002 801 2048
rect 774 1952 777 1998
rect 814 1932 817 2108
rect 848 2103 850 2107
rect 854 2103 857 2107
rect 861 2103 864 2107
rect 870 2072 873 2138
rect 886 2082 889 2148
rect 942 2132 945 2398
rect 950 2362 953 2368
rect 966 2352 969 2458
rect 978 2448 985 2451
rect 982 2392 985 2448
rect 1006 2392 1009 2488
rect 1014 2472 1017 2478
rect 1038 2472 1041 2478
rect 1034 2458 1038 2461
rect 1014 2402 1017 2458
rect 1054 2442 1057 2538
rect 1062 2532 1065 2538
rect 1126 2532 1129 2538
rect 1074 2518 1078 2521
rect 1094 2512 1097 2528
rect 1062 2492 1065 2508
rect 1118 2492 1121 2518
rect 1094 2482 1097 2488
rect 1106 2478 1118 2481
rect 1070 2391 1073 2458
rect 1066 2388 1073 2391
rect 1030 2362 1033 2378
rect 1070 2352 1073 2388
rect 994 2348 998 2351
rect 974 2322 977 2328
rect 1022 2292 1025 2298
rect 1014 2282 1017 2288
rect 978 2268 982 2271
rect 950 2262 953 2268
rect 958 2262 961 2268
rect 970 2258 982 2261
rect 990 2222 993 2278
rect 1002 2258 1006 2261
rect 1030 2242 1033 2348
rect 1046 2322 1049 2338
rect 1038 2281 1041 2318
rect 1038 2278 1046 2281
rect 1062 2262 1065 2268
rect 1070 2262 1073 2278
rect 1078 2272 1081 2358
rect 1086 2262 1089 2468
rect 1110 2442 1113 2468
rect 1118 2452 1121 2458
rect 1126 2442 1129 2518
rect 1142 2472 1145 2618
rect 1150 2552 1153 2568
rect 1166 2562 1169 2688
rect 1222 2672 1225 2678
rect 1238 2662 1241 2668
rect 1290 2658 1294 2661
rect 1302 2652 1305 2728
rect 1310 2682 1313 2718
rect 1182 2561 1185 2638
rect 1222 2592 1225 2648
rect 1270 2631 1273 2650
rect 1294 2612 1297 2638
rect 1182 2558 1193 2561
rect 1182 2542 1185 2548
rect 1190 2542 1193 2558
rect 1206 2552 1209 2568
rect 1246 2552 1249 2598
rect 1274 2558 1278 2561
rect 1158 2522 1161 2538
rect 1198 2522 1201 2538
rect 1222 2531 1225 2548
rect 1218 2528 1225 2531
rect 1230 2542 1233 2548
rect 1262 2542 1265 2548
rect 1294 2542 1297 2608
rect 1242 2538 1246 2541
rect 1230 2532 1233 2538
rect 1150 2482 1153 2518
rect 1166 2482 1169 2518
rect 1230 2508 1238 2511
rect 1230 2492 1233 2508
rect 1218 2488 1222 2491
rect 1254 2482 1257 2538
rect 1270 2532 1273 2538
rect 1286 2512 1289 2518
rect 1162 2468 1166 2471
rect 1146 2458 1150 2461
rect 1134 2392 1137 2458
rect 1142 2332 1145 2418
rect 1174 2412 1177 2458
rect 1182 2432 1185 2478
rect 1206 2472 1209 2478
rect 1202 2458 1206 2461
rect 1206 2442 1209 2448
rect 1222 2432 1225 2448
rect 1230 2442 1233 2448
rect 1190 2360 1193 2379
rect 1202 2348 1206 2351
rect 1078 2252 1081 2258
rect 1094 2251 1097 2298
rect 1102 2282 1105 2288
rect 1110 2272 1113 2288
rect 1158 2281 1161 2338
rect 1190 2292 1193 2318
rect 1222 2292 1225 2408
rect 1246 2342 1249 2478
rect 1270 2442 1273 2468
rect 1278 2412 1281 2458
rect 1286 2422 1289 2468
rect 1254 2392 1257 2398
rect 1270 2352 1273 2358
rect 1294 2352 1297 2398
rect 1310 2362 1313 2458
rect 1318 2442 1321 2738
rect 1334 2652 1337 2658
rect 1342 2572 1345 2718
rect 1350 2702 1353 2738
rect 1422 2712 1425 2748
rect 1438 2742 1441 2748
rect 1390 2672 1393 2678
rect 1406 2672 1409 2678
rect 1358 2622 1361 2650
rect 1406 2621 1409 2668
rect 1446 2662 1449 2668
rect 1398 2618 1409 2621
rect 1360 2603 1362 2607
rect 1366 2603 1369 2607
rect 1373 2603 1376 2607
rect 1350 2560 1353 2579
rect 1382 2552 1385 2558
rect 1342 2492 1345 2518
rect 1360 2403 1362 2407
rect 1366 2403 1369 2407
rect 1373 2403 1376 2407
rect 1326 2392 1329 2398
rect 1382 2362 1385 2538
rect 1398 2532 1401 2618
rect 1398 2511 1401 2528
rect 1390 2508 1401 2511
rect 1310 2352 1313 2358
rect 1170 2288 1174 2291
rect 1158 2278 1169 2281
rect 1118 2272 1121 2278
rect 1150 2262 1153 2268
rect 1106 2258 1110 2261
rect 1086 2248 1097 2251
rect 990 2202 993 2218
rect 1086 2192 1089 2248
rect 1134 2242 1137 2258
rect 990 2160 993 2179
rect 1126 2172 1129 2218
rect 1134 2192 1137 2228
rect 1010 2148 1014 2151
rect 958 2142 961 2148
rect 1102 2142 1105 2168
rect 1130 2158 1134 2161
rect 1110 2152 1113 2158
rect 1126 2142 1129 2148
rect 1150 2142 1153 2158
rect 1034 2138 1038 2141
rect 918 2062 921 2078
rect 890 2058 894 2061
rect 742 1872 745 1928
rect 614 1858 625 1861
rect 634 1858 638 1861
rect 454 1792 457 1848
rect 462 1842 465 1858
rect 494 1852 497 1858
rect 598 1852 601 1858
rect 486 1832 489 1848
rect 470 1762 473 1798
rect 458 1748 462 1751
rect 474 1748 478 1751
rect 486 1742 489 1818
rect 494 1752 497 1848
rect 526 1812 529 1848
rect 502 1752 505 1768
rect 518 1762 521 1778
rect 526 1742 529 1768
rect 550 1762 553 1808
rect 558 1762 561 1848
rect 578 1838 582 1841
rect 566 1832 569 1838
rect 614 1822 617 1848
rect 570 1778 574 1781
rect 570 1768 574 1771
rect 562 1758 577 1761
rect 546 1748 550 1751
rect 562 1748 566 1751
rect 534 1742 537 1748
rect 418 1738 422 1741
rect 434 1738 441 1741
rect 406 1692 409 1698
rect 394 1678 401 1681
rect 382 1578 393 1581
rect 382 1562 385 1568
rect 390 1562 393 1578
rect 398 1542 401 1678
rect 414 1552 417 1738
rect 426 1728 430 1731
rect 438 1692 441 1738
rect 446 1702 449 1738
rect 486 1722 489 1738
rect 486 1692 489 1708
rect 494 1702 497 1738
rect 510 1701 513 1738
rect 526 1732 529 1738
rect 574 1722 577 1758
rect 502 1698 513 1701
rect 486 1682 489 1688
rect 502 1672 505 1698
rect 582 1692 585 1808
rect 622 1762 625 1858
rect 654 1852 657 1868
rect 742 1862 745 1868
rect 722 1858 729 1861
rect 674 1848 678 1851
rect 646 1832 649 1848
rect 630 1792 633 1798
rect 642 1768 646 1771
rect 654 1762 657 1838
rect 686 1792 689 1858
rect 718 1852 721 1858
rect 702 1832 705 1848
rect 590 1752 593 1758
rect 622 1722 625 1758
rect 634 1748 638 1751
rect 654 1742 657 1748
rect 662 1732 665 1758
rect 674 1748 678 1751
rect 686 1742 689 1768
rect 694 1752 697 1768
rect 674 1738 678 1741
rect 598 1672 601 1698
rect 606 1682 609 1718
rect 618 1668 622 1671
rect 442 1658 446 1661
rect 534 1631 537 1650
rect 454 1592 457 1598
rect 510 1592 513 1618
rect 470 1582 473 1588
rect 490 1558 494 1561
rect 438 1552 441 1558
rect 510 1548 518 1551
rect 462 1542 465 1548
rect 434 1538 438 1541
rect 382 1512 385 1518
rect 390 1492 393 1518
rect 406 1502 409 1538
rect 446 1532 449 1538
rect 370 1478 377 1481
rect 382 1482 385 1488
rect 390 1472 393 1488
rect 398 1462 401 1478
rect 414 1472 417 1528
rect 422 1482 425 1518
rect 426 1468 430 1471
rect 402 1448 406 1451
rect 414 1432 417 1468
rect 430 1442 433 1448
rect 344 1403 346 1407
rect 350 1403 353 1407
rect 357 1403 360 1407
rect 374 1392 377 1418
rect 438 1412 441 1498
rect 454 1482 457 1538
rect 494 1522 497 1548
rect 510 1512 513 1548
rect 522 1538 526 1541
rect 510 1492 513 1508
rect 526 1492 529 1538
rect 542 1492 545 1658
rect 574 1652 577 1658
rect 574 1622 577 1648
rect 590 1632 593 1668
rect 602 1658 606 1661
rect 598 1612 601 1658
rect 630 1652 633 1718
rect 678 1692 681 1728
rect 638 1662 641 1688
rect 686 1672 689 1738
rect 694 1722 697 1748
rect 710 1702 713 1718
rect 646 1642 649 1668
rect 662 1662 665 1668
rect 710 1652 713 1658
rect 550 1562 553 1588
rect 570 1568 574 1571
rect 558 1562 561 1568
rect 590 1562 593 1578
rect 582 1552 585 1558
rect 606 1552 609 1628
rect 574 1542 577 1548
rect 590 1542 593 1548
rect 606 1542 609 1548
rect 614 1542 617 1598
rect 646 1572 649 1638
rect 654 1552 657 1648
rect 682 1638 686 1641
rect 670 1582 673 1618
rect 718 1612 721 1668
rect 726 1662 729 1858
rect 762 1848 766 1851
rect 734 1822 737 1848
rect 734 1712 737 1818
rect 750 1742 753 1748
rect 758 1742 761 1758
rect 766 1742 769 1748
rect 750 1722 753 1738
rect 762 1728 766 1731
rect 742 1701 745 1718
rect 734 1698 745 1701
rect 694 1582 697 1588
rect 674 1568 678 1571
rect 698 1568 702 1571
rect 622 1522 625 1548
rect 638 1532 641 1538
rect 446 1432 449 1468
rect 454 1461 457 1478
rect 462 1472 465 1488
rect 522 1478 526 1481
rect 478 1472 481 1478
rect 534 1472 537 1478
rect 490 1468 494 1471
rect 454 1458 465 1461
rect 334 1352 337 1378
rect 350 1360 353 1379
rect 334 1332 337 1348
rect 382 1342 385 1398
rect 398 1322 401 1328
rect 446 1302 449 1428
rect 382 1272 385 1278
rect 398 1272 401 1278
rect 342 1262 345 1268
rect 454 1262 457 1438
rect 446 1222 449 1248
rect 454 1222 457 1258
rect 344 1203 346 1207
rect 350 1203 353 1207
rect 357 1203 360 1207
rect 342 1142 345 1148
rect 278 1092 281 1098
rect 246 1078 257 1081
rect 230 1072 233 1078
rect 50 1058 54 1061
rect 30 1048 41 1051
rect 30 952 33 1048
rect 70 960 73 1048
rect 118 982 121 1068
rect 230 1062 233 1068
rect 246 1062 249 1068
rect 254 1061 257 1078
rect 254 1058 262 1061
rect 174 1031 177 1058
rect 254 1052 257 1058
rect 14 852 17 918
rect 30 752 33 948
rect 46 922 49 958
rect 102 952 105 978
rect 102 932 105 938
rect 214 932 217 1018
rect 238 992 241 1018
rect 238 972 241 978
rect 262 962 265 1018
rect 286 962 289 1138
rect 310 1122 313 1128
rect 318 1102 321 1128
rect 294 1042 297 1058
rect 302 1052 305 1058
rect 310 1052 313 1088
rect 326 1082 329 1108
rect 334 1092 337 1138
rect 342 1122 345 1138
rect 358 1092 361 1138
rect 322 1058 326 1061
rect 322 1048 326 1051
rect 310 1042 313 1048
rect 302 982 305 1018
rect 344 1003 346 1007
rect 350 1003 353 1007
rect 357 1003 360 1007
rect 374 992 377 1218
rect 462 1192 465 1458
rect 470 1452 473 1458
rect 486 1452 489 1458
rect 502 1372 505 1468
rect 518 1392 521 1408
rect 490 1368 494 1371
rect 502 1332 505 1368
rect 534 1362 537 1458
rect 550 1402 553 1518
rect 614 1472 617 1478
rect 630 1472 633 1478
rect 566 1422 569 1448
rect 574 1442 577 1458
rect 598 1392 601 1398
rect 658 1388 662 1391
rect 554 1368 558 1371
rect 578 1368 582 1371
rect 510 1342 513 1348
rect 526 1342 529 1348
rect 470 1282 473 1288
rect 502 1272 505 1278
rect 482 1268 486 1271
rect 498 1258 502 1261
rect 478 1172 481 1218
rect 510 1192 513 1328
rect 534 1312 537 1358
rect 542 1352 545 1358
rect 542 1332 545 1338
rect 562 1328 566 1331
rect 534 1272 537 1298
rect 542 1292 545 1318
rect 582 1312 585 1348
rect 590 1342 593 1348
rect 574 1308 582 1311
rect 518 1252 521 1268
rect 534 1252 537 1268
rect 522 1168 526 1171
rect 538 1168 542 1171
rect 430 1162 433 1168
rect 502 1162 505 1168
rect 478 1152 481 1158
rect 510 1152 513 1158
rect 426 1148 430 1151
rect 442 1148 446 1151
rect 538 1148 542 1151
rect 454 1142 457 1148
rect 494 1142 497 1148
rect 558 1142 561 1268
rect 566 1262 569 1268
rect 442 1138 446 1141
rect 422 1112 425 1138
rect 454 1122 457 1138
rect 470 1122 473 1138
rect 550 1132 553 1138
rect 462 1102 465 1118
rect 438 1072 441 1078
rect 454 1072 457 1088
rect 398 1031 401 1058
rect 422 992 425 998
rect 326 962 329 968
rect 290 958 294 961
rect 390 952 393 978
rect 314 948 318 951
rect 338 948 342 951
rect 222 938 230 941
rect 266 938 270 941
rect 306 938 310 941
rect 118 902 121 928
rect 198 902 201 918
rect 86 882 89 888
rect 214 882 217 928
rect 222 892 225 938
rect 238 892 241 908
rect 70 862 73 868
rect 126 831 129 858
rect 182 842 185 878
rect 170 818 174 821
rect 186 778 190 781
rect 198 772 201 868
rect 226 848 230 851
rect 54 762 57 768
rect 74 748 78 751
rect 98 738 102 741
rect 78 732 81 738
rect 126 731 129 768
rect 134 742 137 748
rect 158 742 161 768
rect 178 758 185 761
rect 146 738 150 741
rect 126 728 134 731
rect 146 728 150 731
rect 14 652 17 718
rect 86 702 89 718
rect 70 672 73 698
rect 86 682 89 688
rect 166 682 169 748
rect 170 678 174 681
rect 182 662 185 758
rect 190 682 193 748
rect 198 742 201 768
rect 206 752 209 778
rect 214 742 217 748
rect 254 742 257 818
rect 262 752 265 838
rect 270 752 273 918
rect 278 792 281 868
rect 286 761 289 918
rect 310 882 313 888
rect 334 882 337 888
rect 298 868 302 871
rect 342 862 345 948
rect 322 858 326 861
rect 302 782 305 818
rect 314 768 318 771
rect 286 758 294 761
rect 302 752 305 758
rect 282 748 286 751
rect 234 738 238 741
rect 242 728 246 731
rect 218 718 222 721
rect 230 712 233 728
rect 238 701 241 728
rect 262 722 265 748
rect 230 698 241 701
rect 202 678 206 681
rect 202 668 206 671
rect 174 658 182 661
rect 202 658 206 661
rect 14 562 17 648
rect 126 631 129 658
rect 174 591 177 658
rect 170 588 177 591
rect 38 560 41 561
rect 14 392 17 528
rect 38 454 41 556
rect 70 552 73 578
rect 206 562 209 578
rect 214 562 217 568
rect 194 548 201 551
rect 182 542 185 548
rect 70 522 73 538
rect 86 522 89 528
rect 198 492 201 548
rect 222 522 225 678
rect 230 552 233 698
rect 238 682 241 688
rect 246 672 249 718
rect 242 668 246 671
rect 254 662 257 698
rect 270 692 273 738
rect 278 732 281 748
rect 294 692 297 748
rect 278 672 281 678
rect 246 562 249 568
rect 230 542 233 548
rect 206 502 209 518
rect 214 512 217 518
rect 222 492 225 518
rect 238 492 241 538
rect 170 488 174 491
rect 70 472 73 488
rect 86 472 89 478
rect 230 472 233 488
rect 246 482 249 518
rect 254 512 257 658
rect 178 468 182 471
rect 262 462 265 668
rect 278 592 281 668
rect 278 552 281 558
rect 286 552 289 558
rect 302 552 305 748
rect 310 662 313 688
rect 318 682 321 728
rect 326 692 329 858
rect 366 822 369 878
rect 382 862 385 878
rect 390 862 393 938
rect 430 932 433 938
rect 406 922 409 928
rect 438 892 441 1028
rect 454 992 457 1038
rect 486 1022 489 1118
rect 506 1048 510 1051
rect 446 932 449 968
rect 494 962 497 968
rect 466 958 470 961
rect 474 948 478 951
rect 454 942 457 948
rect 534 942 537 1018
rect 550 992 553 1128
rect 558 1122 561 1138
rect 574 1071 577 1308
rect 582 1272 585 1288
rect 590 1282 593 1298
rect 582 1202 585 1238
rect 582 1152 585 1198
rect 598 1192 601 1348
rect 626 1338 630 1341
rect 646 1262 649 1378
rect 670 1342 673 1488
rect 678 1372 681 1568
rect 686 1362 689 1558
rect 718 1552 721 1568
rect 698 1548 702 1551
rect 710 1492 713 1528
rect 718 1512 721 1538
rect 726 1512 729 1658
rect 734 1652 737 1698
rect 742 1682 745 1688
rect 746 1668 750 1671
rect 758 1662 761 1718
rect 766 1672 769 1688
rect 774 1682 777 1908
rect 806 1892 809 1908
rect 814 1872 817 1918
rect 830 1911 833 1938
rect 862 1922 865 2038
rect 878 2002 881 2058
rect 906 2038 910 2041
rect 878 1962 881 1988
rect 830 1908 841 1911
rect 838 1891 841 1908
rect 848 1903 850 1907
rect 854 1903 857 1907
rect 861 1903 864 1907
rect 838 1888 846 1891
rect 822 1872 825 1878
rect 838 1872 841 1878
rect 786 1868 790 1871
rect 786 1858 790 1861
rect 794 1848 798 1851
rect 850 1848 854 1851
rect 782 1742 785 1818
rect 806 1792 809 1828
rect 798 1772 801 1788
rect 814 1772 817 1838
rect 822 1802 825 1848
rect 862 1781 865 1868
rect 894 1862 897 2028
rect 914 1958 918 1961
rect 926 1952 929 2048
rect 942 2042 945 2108
rect 950 2062 953 2088
rect 958 2052 961 2118
rect 1046 2082 1049 2138
rect 1130 2088 1134 2091
rect 1142 2082 1145 2128
rect 1158 2092 1161 2238
rect 1166 2152 1169 2278
rect 1174 2272 1177 2278
rect 1198 2252 1201 2258
rect 1182 2182 1185 2248
rect 1202 2238 1206 2241
rect 1230 2192 1233 2328
rect 1246 2272 1249 2338
rect 1270 2332 1273 2348
rect 1334 2342 1337 2348
rect 1306 2338 1310 2341
rect 1322 2338 1326 2341
rect 1278 2312 1281 2338
rect 1286 2332 1289 2338
rect 1338 2328 1342 2331
rect 1246 2251 1249 2268
rect 1238 2248 1249 2251
rect 1302 2262 1305 2278
rect 1318 2272 1321 2278
rect 1366 2262 1369 2348
rect 1382 2332 1385 2338
rect 1374 2322 1377 2328
rect 1382 2312 1385 2328
rect 1374 2301 1377 2308
rect 1390 2302 1393 2508
rect 1402 2488 1406 2491
rect 1442 2468 1446 2471
rect 1406 2462 1409 2468
rect 1434 2458 1438 2461
rect 1422 2432 1425 2438
rect 1470 2412 1473 2748
rect 1478 2742 1481 2758
rect 1490 2738 1494 2741
rect 1486 2701 1489 2718
rect 1478 2698 1489 2701
rect 1478 2602 1481 2698
rect 1490 2688 1494 2691
rect 1502 2582 1505 2818
rect 1518 2792 1521 2808
rect 1510 2732 1513 2748
rect 1526 2722 1529 2818
rect 1534 2711 1537 2908
rect 1558 2881 1561 2938
rect 1566 2922 1569 2948
rect 1590 2942 1593 2948
rect 1630 2942 1633 2998
rect 1646 2942 1649 3078
rect 1654 2942 1657 3148
rect 1690 3138 1694 3141
rect 1662 3082 1665 3118
rect 1674 3088 1678 3091
rect 1694 3072 1697 3098
rect 1702 3072 1705 3288
rect 1790 3282 1793 3288
rect 1710 3212 1713 3218
rect 1722 3188 1726 3191
rect 1718 3168 1726 3171
rect 1710 3152 1713 3158
rect 1718 3092 1721 3168
rect 1734 3122 1737 3148
rect 1750 3112 1753 3158
rect 1766 3142 1769 3208
rect 1806 3202 1809 3268
rect 1838 3222 1841 3250
rect 1846 3192 1849 3258
rect 1870 3252 1873 3288
rect 2006 3282 2009 3388
rect 2054 3352 2057 3408
rect 2086 3392 2089 3418
rect 2014 3312 2017 3318
rect 1906 3268 1910 3271
rect 1890 3248 1894 3251
rect 1790 3162 1793 3168
rect 1798 3162 1801 3168
rect 1814 3162 1817 3168
rect 1778 3138 1782 3141
rect 1798 3132 1801 3138
rect 1734 3072 1737 3078
rect 1758 3072 1761 3108
rect 1714 3068 1718 3071
rect 1662 2992 1665 3068
rect 1670 3052 1673 3068
rect 1690 3058 1694 3061
rect 1674 3048 1681 3051
rect 1550 2878 1561 2881
rect 1606 2882 1609 2938
rect 1638 2902 1641 2918
rect 1550 2742 1553 2878
rect 1622 2862 1625 2868
rect 1662 2862 1665 2988
rect 1670 2962 1673 2978
rect 1678 2962 1681 3048
rect 1718 2992 1721 3018
rect 1670 2922 1673 2928
rect 1526 2708 1537 2711
rect 1526 2682 1529 2708
rect 1534 2682 1537 2688
rect 1558 2672 1561 2748
rect 1614 2742 1617 2758
rect 1654 2752 1657 2858
rect 1670 2822 1673 2848
rect 1678 2802 1681 2958
rect 1694 2952 1697 2958
rect 1694 2901 1697 2938
rect 1694 2898 1702 2901
rect 1710 2892 1713 2968
rect 1718 2952 1721 2958
rect 1726 2952 1729 2958
rect 1698 2868 1702 2871
rect 1722 2868 1726 2871
rect 1734 2871 1737 3058
rect 1742 3052 1745 3058
rect 1758 3052 1761 3068
rect 1782 3052 1785 3128
rect 1790 3052 1793 3118
rect 1822 3102 1825 3138
rect 1830 3062 1833 3188
rect 1866 3158 1870 3161
rect 1886 3152 1889 3198
rect 1902 3162 1905 3218
rect 1926 3202 1929 3218
rect 2022 3202 2025 3268
rect 2054 3262 2057 3348
rect 2094 3332 2097 3488
rect 2142 3472 2145 3488
rect 2150 3452 2153 3458
rect 2166 3442 2169 3448
rect 2182 3412 2185 3478
rect 2202 3468 2206 3471
rect 2222 3462 2225 3548
rect 2262 3542 2265 3568
rect 2370 3558 2374 3561
rect 2402 3558 2406 3561
rect 2430 3552 2433 3588
rect 2450 3568 2454 3571
rect 2478 3562 2481 3568
rect 2466 3558 2470 3561
rect 2542 3560 2545 3579
rect 2702 3562 2705 3588
rect 2446 3552 2449 3558
rect 2506 3548 2510 3551
rect 2422 3542 2425 3548
rect 2386 3538 2390 3541
rect 2278 3532 2281 3538
rect 2230 3492 2233 3508
rect 2246 3492 2249 3508
rect 2238 3472 2241 3478
rect 2254 3472 2257 3488
rect 2262 3472 2265 3528
rect 2358 3522 2361 3538
rect 2430 3522 2433 3548
rect 2350 3518 2358 3521
rect 2278 3492 2281 3508
rect 2270 3482 2273 3488
rect 2350 3482 2353 3518
rect 2438 3512 2441 3538
rect 2462 3512 2465 3548
rect 2630 3542 2633 3548
rect 2702 3542 2705 3548
rect 2750 3542 2753 3558
rect 2474 3538 2478 3541
rect 2494 3532 2497 3538
rect 2574 3532 2577 3538
rect 2438 3482 2441 3498
rect 2526 3482 2529 3508
rect 2590 3502 2593 3528
rect 2670 3512 2673 3518
rect 2302 3472 2305 3478
rect 2194 3458 2198 3461
rect 2266 3458 2270 3461
rect 2214 3452 2217 3458
rect 2190 3392 2193 3448
rect 2142 3360 2145 3379
rect 2254 3352 2257 3458
rect 2306 3418 2310 3421
rect 2178 3348 2182 3351
rect 2150 3341 2153 3348
rect 2142 3338 2153 3341
rect 2110 3332 2113 3338
rect 2094 3282 2097 3328
rect 2070 3222 2073 3248
rect 2102 3202 2105 3218
rect 2038 3192 2041 3198
rect 1842 3148 1846 3151
rect 1926 3142 1929 3148
rect 1934 3142 1937 3168
rect 1958 3152 1961 3158
rect 1966 3142 1969 3168
rect 1998 3162 2001 3168
rect 2110 3162 2113 3168
rect 2066 3158 2070 3161
rect 2082 3158 2086 3161
rect 1978 3148 1982 3151
rect 1990 3142 1993 3148
rect 1890 3138 1894 3141
rect 1838 3132 1841 3138
rect 1880 3103 1882 3107
rect 1886 3103 1889 3107
rect 1893 3103 1896 3107
rect 1870 3082 1873 3088
rect 1766 3032 1769 3038
rect 1790 3002 1793 3018
rect 1830 2992 1833 3058
rect 1886 3042 1889 3068
rect 1782 2952 1785 2988
rect 1870 2960 1873 2979
rect 1838 2932 1841 2938
rect 1742 2912 1745 2918
rect 1822 2902 1825 2928
rect 1880 2903 1882 2907
rect 1886 2903 1889 2907
rect 1893 2903 1896 2907
rect 1854 2882 1857 2898
rect 1746 2878 1750 2881
rect 1734 2868 1745 2871
rect 1662 2762 1665 2788
rect 1694 2752 1697 2858
rect 1734 2792 1737 2858
rect 1742 2832 1745 2868
rect 1758 2812 1761 2858
rect 1766 2802 1769 2858
rect 1854 2852 1857 2878
rect 1710 2772 1713 2778
rect 1730 2768 1734 2771
rect 1758 2762 1761 2798
rect 1726 2752 1729 2758
rect 1682 2748 1686 2751
rect 1746 2748 1750 2751
rect 1566 2682 1569 2688
rect 1574 2672 1577 2678
rect 1586 2668 1590 2671
rect 1554 2658 1558 2661
rect 1510 2652 1513 2658
rect 1518 2582 1521 2618
rect 1542 2572 1545 2598
rect 1550 2592 1553 2618
rect 1582 2612 1585 2658
rect 1598 2632 1601 2728
rect 1686 2722 1689 2748
rect 1706 2738 1710 2741
rect 1694 2732 1697 2738
rect 1718 2711 1721 2748
rect 1774 2742 1777 2818
rect 1782 2762 1785 2768
rect 1798 2742 1801 2818
rect 1854 2802 1857 2848
rect 1846 2792 1849 2798
rect 1822 2762 1825 2788
rect 1718 2708 1726 2711
rect 1618 2668 1622 2671
rect 1598 2592 1601 2618
rect 1614 2602 1617 2658
rect 1630 2652 1633 2698
rect 1642 2688 1646 2691
rect 1722 2688 1726 2691
rect 1654 2662 1657 2668
rect 1638 2652 1641 2658
rect 1662 2632 1665 2668
rect 1670 2652 1673 2688
rect 1758 2682 1761 2688
rect 1678 2672 1681 2678
rect 1694 2672 1697 2678
rect 1714 2668 1718 2671
rect 1686 2662 1689 2668
rect 1702 2652 1705 2658
rect 1726 2612 1729 2678
rect 1774 2672 1777 2738
rect 1782 2692 1785 2708
rect 1790 2702 1793 2718
rect 1798 2672 1801 2738
rect 1806 2732 1809 2738
rect 1814 2681 1817 2728
rect 1806 2678 1817 2681
rect 1806 2672 1809 2678
rect 1838 2672 1841 2788
rect 1846 2742 1849 2748
rect 1854 2692 1857 2758
rect 1862 2712 1865 2728
rect 1738 2668 1742 2671
rect 1734 2632 1737 2648
rect 1582 2562 1585 2588
rect 1750 2582 1753 2668
rect 1514 2558 1518 2561
rect 1530 2558 1537 2561
rect 1510 2542 1513 2548
rect 1498 2538 1502 2541
rect 1502 2472 1505 2518
rect 1518 2472 1521 2478
rect 1526 2462 1529 2488
rect 1534 2442 1537 2558
rect 1550 2542 1553 2548
rect 1542 2492 1545 2528
rect 1558 2492 1561 2558
rect 1758 2552 1761 2658
rect 1766 2562 1769 2618
rect 1578 2548 1582 2551
rect 1766 2542 1769 2548
rect 1774 2542 1777 2548
rect 1542 2452 1545 2458
rect 1498 2418 1502 2421
rect 1550 2412 1553 2468
rect 1558 2442 1561 2448
rect 1574 2382 1577 2468
rect 1582 2422 1585 2468
rect 1510 2360 1513 2379
rect 1418 2348 1422 2351
rect 1478 2332 1481 2338
rect 1462 2302 1465 2328
rect 1374 2298 1385 2301
rect 1218 2188 1222 2191
rect 1190 2142 1193 2148
rect 1170 2138 1174 2141
rect 1202 2138 1206 2141
rect 1190 2092 1193 2138
rect 1198 2092 1201 2108
rect 1030 2072 1033 2078
rect 1046 2072 1049 2078
rect 982 2052 985 2058
rect 934 1952 937 1968
rect 902 1902 905 1918
rect 942 1912 945 2038
rect 950 2022 953 2028
rect 950 1992 953 1998
rect 958 1972 961 2048
rect 998 2031 1001 2050
rect 1014 1992 1017 2008
rect 1030 1992 1033 1998
rect 1070 1992 1073 1998
rect 1126 1992 1129 2078
rect 1214 2072 1217 2178
rect 1230 2102 1233 2188
rect 1238 2112 1241 2248
rect 1214 2062 1217 2068
rect 1078 1972 1081 1988
rect 1102 1972 1105 1978
rect 1134 1972 1137 1978
rect 1066 1968 1070 1971
rect 994 1958 998 1961
rect 1054 1952 1057 1958
rect 986 1948 990 1951
rect 1006 1948 1014 1951
rect 902 1862 905 1898
rect 918 1852 921 1878
rect 926 1872 929 1878
rect 934 1872 937 1878
rect 870 1792 873 1848
rect 898 1838 902 1841
rect 910 1832 913 1848
rect 902 1802 905 1818
rect 942 1812 945 1858
rect 950 1852 953 1918
rect 958 1902 961 1928
rect 962 1868 966 1871
rect 962 1848 966 1851
rect 974 1792 977 1918
rect 1006 1902 1009 1948
rect 1018 1938 1022 1941
rect 986 1858 990 1861
rect 998 1852 1001 1868
rect 986 1838 990 1841
rect 998 1832 1001 1848
rect 990 1782 993 1818
rect 862 1778 873 1781
rect 798 1762 801 1768
rect 790 1752 793 1758
rect 790 1732 793 1738
rect 782 1728 790 1731
rect 782 1672 785 1728
rect 770 1658 774 1661
rect 746 1648 750 1651
rect 758 1592 761 1608
rect 750 1562 753 1578
rect 738 1548 742 1551
rect 790 1542 793 1678
rect 806 1672 809 1748
rect 814 1712 817 1768
rect 822 1692 825 1758
rect 846 1752 849 1758
rect 854 1752 857 1768
rect 834 1748 838 1751
rect 830 1722 833 1738
rect 802 1658 806 1661
rect 822 1582 825 1648
rect 830 1592 833 1708
rect 848 1703 850 1707
rect 854 1703 857 1707
rect 861 1703 864 1707
rect 870 1702 873 1778
rect 918 1752 921 1778
rect 986 1768 990 1771
rect 998 1752 1001 1758
rect 882 1748 886 1751
rect 978 1748 982 1751
rect 914 1738 918 1741
rect 878 1692 881 1718
rect 842 1668 846 1671
rect 838 1632 841 1658
rect 818 1548 822 1551
rect 746 1528 750 1531
rect 758 1528 766 1531
rect 726 1492 729 1498
rect 742 1452 745 1468
rect 750 1462 753 1518
rect 726 1422 729 1438
rect 726 1382 729 1418
rect 714 1368 718 1371
rect 734 1362 737 1418
rect 742 1401 745 1448
rect 758 1432 761 1528
rect 766 1492 769 1508
rect 790 1492 793 1538
rect 802 1528 806 1531
rect 834 1528 838 1531
rect 862 1522 865 1548
rect 798 1512 801 1518
rect 848 1503 850 1507
rect 854 1503 857 1507
rect 861 1503 864 1507
rect 766 1482 769 1488
rect 838 1472 841 1488
rect 870 1472 873 1568
rect 886 1542 889 1738
rect 910 1732 913 1738
rect 902 1722 905 1728
rect 910 1671 913 1728
rect 926 1722 929 1738
rect 922 1688 926 1691
rect 934 1682 937 1748
rect 950 1742 953 1748
rect 942 1732 945 1738
rect 998 1732 1001 1738
rect 990 1722 993 1728
rect 950 1692 953 1708
rect 942 1682 945 1688
rect 966 1682 969 1718
rect 1006 1682 1009 1758
rect 1014 1692 1017 1928
rect 1030 1862 1033 1868
rect 1038 1752 1041 1918
rect 1046 1872 1049 1948
rect 1054 1882 1057 1948
rect 1054 1872 1057 1878
rect 1046 1852 1049 1868
rect 1062 1862 1065 1968
rect 1126 1962 1129 1968
rect 1114 1958 1118 1961
rect 1074 1948 1078 1951
rect 1094 1942 1097 1948
rect 1118 1942 1121 1958
rect 1126 1952 1129 1958
rect 1142 1952 1145 2048
rect 1022 1692 1025 1748
rect 1058 1738 1062 1741
rect 1030 1722 1033 1738
rect 906 1668 913 1671
rect 926 1662 929 1678
rect 934 1662 937 1668
rect 1030 1662 1033 1668
rect 1038 1662 1041 1728
rect 1070 1722 1073 1918
rect 1078 1882 1081 1888
rect 1078 1862 1081 1878
rect 1098 1868 1102 1871
rect 1102 1832 1105 1858
rect 1118 1852 1121 1928
rect 1126 1872 1129 1948
rect 1150 1932 1153 2058
rect 1174 2042 1177 2048
rect 1158 2002 1161 2038
rect 1182 2002 1185 2058
rect 1206 2042 1209 2048
rect 1194 2038 1198 2041
rect 1182 1992 1185 1998
rect 1166 1982 1169 1988
rect 1190 1972 1193 2038
rect 1158 1962 1161 1968
rect 1166 1952 1169 1968
rect 1198 1962 1201 2018
rect 1214 1962 1217 1988
rect 1142 1872 1145 1918
rect 1158 1872 1161 1948
rect 1174 1932 1177 1958
rect 1222 1942 1225 2078
rect 1238 2062 1241 2078
rect 1246 2072 1249 2238
rect 1302 2221 1305 2258
rect 1350 2231 1353 2250
rect 1294 2218 1305 2221
rect 1254 2142 1257 2148
rect 1294 2132 1297 2218
rect 1360 2203 1362 2207
rect 1366 2203 1369 2207
rect 1373 2203 1376 2207
rect 1382 2192 1385 2298
rect 1518 2292 1521 2328
rect 1466 2288 1470 2291
rect 1406 2272 1409 2288
rect 1414 2282 1417 2288
rect 1422 2262 1425 2268
rect 1430 2251 1433 2288
rect 1502 2272 1505 2278
rect 1450 2268 1454 2271
rect 1514 2268 1518 2271
rect 1522 2268 1533 2271
rect 1494 2262 1497 2268
rect 1426 2248 1433 2251
rect 1358 2162 1361 2188
rect 1438 2182 1441 2188
rect 1310 2142 1313 2148
rect 1294 2122 1297 2128
rect 1278 2092 1281 2108
rect 1310 2092 1313 2128
rect 1362 2068 1366 2071
rect 1258 2058 1262 2061
rect 1238 2032 1241 2058
rect 1294 2022 1297 2058
rect 1230 1972 1233 2018
rect 1254 2012 1257 2018
rect 1322 1948 1326 1951
rect 1186 1938 1190 1941
rect 1206 1882 1209 1908
rect 1222 1892 1225 1938
rect 1230 1892 1233 1928
rect 1214 1882 1217 1888
rect 1194 1878 1198 1881
rect 1114 1848 1118 1851
rect 1078 1792 1081 1808
rect 906 1658 910 1661
rect 994 1658 998 1661
rect 894 1562 897 1658
rect 914 1588 918 1591
rect 946 1588 950 1591
rect 958 1552 961 1598
rect 966 1592 969 1658
rect 982 1652 985 1658
rect 982 1602 985 1618
rect 982 1552 985 1568
rect 998 1562 1001 1598
rect 1006 1592 1009 1648
rect 878 1522 881 1538
rect 894 1522 897 1548
rect 878 1512 881 1518
rect 858 1468 862 1471
rect 798 1462 801 1468
rect 814 1462 817 1468
rect 834 1458 838 1461
rect 846 1452 849 1458
rect 806 1442 809 1448
rect 742 1398 750 1401
rect 706 1358 710 1361
rect 750 1352 753 1398
rect 790 1372 793 1438
rect 814 1432 817 1448
rect 798 1412 801 1418
rect 802 1368 806 1371
rect 822 1362 825 1438
rect 854 1432 857 1438
rect 854 1362 857 1408
rect 874 1388 878 1391
rect 894 1382 897 1418
rect 826 1358 830 1361
rect 682 1348 686 1351
rect 778 1348 785 1351
rect 718 1341 721 1348
rect 758 1342 761 1348
rect 718 1338 734 1341
rect 770 1338 774 1341
rect 686 1282 689 1328
rect 694 1302 697 1318
rect 610 1238 614 1241
rect 606 1152 609 1238
rect 686 1192 689 1278
rect 702 1272 705 1278
rect 746 1258 750 1261
rect 734 1231 737 1250
rect 710 1152 713 1178
rect 742 1160 745 1218
rect 590 1132 593 1138
rect 710 1132 713 1138
rect 614 1112 617 1118
rect 694 1092 697 1128
rect 758 1122 761 1338
rect 782 1292 785 1348
rect 826 1348 830 1351
rect 790 1272 793 1318
rect 774 1242 777 1268
rect 798 1142 801 1318
rect 814 1282 817 1348
rect 826 1338 830 1341
rect 894 1332 897 1348
rect 902 1342 905 1528
rect 926 1522 929 1548
rect 958 1532 961 1538
rect 910 1431 913 1518
rect 918 1462 921 1518
rect 934 1462 937 1468
rect 910 1428 921 1431
rect 918 1372 921 1428
rect 942 1402 945 1518
rect 966 1482 969 1498
rect 966 1472 969 1478
rect 974 1472 977 1528
rect 990 1482 993 1538
rect 1014 1522 1017 1538
rect 1002 1488 1006 1491
rect 1006 1472 1009 1478
rect 1014 1472 1017 1508
rect 1022 1492 1025 1578
rect 1038 1552 1041 1658
rect 1046 1562 1049 1718
rect 1094 1692 1097 1728
rect 1110 1692 1113 1848
rect 1142 1832 1145 1858
rect 1222 1852 1225 1858
rect 1178 1848 1182 1851
rect 1158 1732 1161 1818
rect 1222 1762 1225 1788
rect 1226 1748 1230 1751
rect 1174 1722 1177 1738
rect 1206 1692 1209 1708
rect 1054 1682 1057 1688
rect 1070 1682 1073 1688
rect 1118 1672 1121 1678
rect 1182 1672 1185 1678
rect 1110 1662 1113 1668
rect 1090 1658 1094 1661
rect 1142 1652 1145 1658
rect 1158 1642 1161 1648
rect 1174 1632 1177 1668
rect 1198 1652 1201 1688
rect 1206 1662 1209 1668
rect 1190 1632 1193 1638
rect 1110 1562 1113 1608
rect 1082 1558 1086 1561
rect 1046 1552 1049 1558
rect 1054 1552 1057 1558
rect 1126 1542 1129 1628
rect 1170 1618 1174 1621
rect 1134 1562 1137 1618
rect 1158 1592 1161 1598
rect 1198 1591 1201 1648
rect 1214 1642 1217 1738
rect 1238 1712 1241 1868
rect 1246 1852 1249 1858
rect 1262 1852 1265 1938
rect 1278 1872 1281 1928
rect 1318 1892 1321 1918
rect 1270 1842 1273 1868
rect 1294 1862 1297 1878
rect 1282 1848 1289 1851
rect 1286 1792 1289 1848
rect 1302 1832 1305 1868
rect 1326 1832 1329 1878
rect 1334 1872 1337 2068
rect 1390 2062 1393 2118
rect 1406 2101 1409 2128
rect 1406 2098 1417 2101
rect 1406 2082 1409 2088
rect 1360 2003 1362 2007
rect 1366 2003 1369 2007
rect 1373 2003 1376 2007
rect 1354 1988 1358 1991
rect 1390 1922 1393 2058
rect 1398 1942 1401 1948
rect 1406 1942 1409 2018
rect 1414 1992 1417 2098
rect 1422 2092 1425 2098
rect 1422 2072 1425 2088
rect 1422 1991 1425 2018
rect 1430 2002 1433 2018
rect 1438 2012 1441 2168
rect 1446 2162 1449 2258
rect 1478 2232 1481 2248
rect 1518 2202 1521 2218
rect 1526 2192 1529 2248
rect 1458 2148 1462 2151
rect 1458 2138 1462 2141
rect 1446 2132 1449 2138
rect 1470 2082 1473 2158
rect 1494 2152 1497 2158
rect 1510 2142 1513 2158
rect 1486 2122 1489 2138
rect 1494 2132 1497 2138
rect 1466 2078 1470 2081
rect 1446 2062 1449 2068
rect 1462 2062 1465 2068
rect 1470 2062 1473 2068
rect 1422 1988 1433 1991
rect 1430 1962 1433 1988
rect 1446 1952 1449 2058
rect 1458 2048 1462 2051
rect 1470 1992 1473 2038
rect 1478 1972 1481 2118
rect 1518 2112 1521 2138
rect 1510 2101 1513 2108
rect 1510 2098 1521 2101
rect 1486 2072 1489 2078
rect 1494 2062 1497 2098
rect 1518 2092 1521 2098
rect 1534 2082 1537 2088
rect 1502 2062 1505 2068
rect 1510 2042 1513 2068
rect 1542 1992 1545 2378
rect 1562 2358 1566 2361
rect 1562 2348 1566 2351
rect 1574 2342 1577 2358
rect 1590 2352 1593 2498
rect 1630 2492 1633 2538
rect 1646 2522 1649 2528
rect 1638 2498 1646 2501
rect 1638 2492 1641 2498
rect 1650 2468 1654 2471
rect 1662 2462 1665 2508
rect 1602 2358 1606 2361
rect 1550 2252 1553 2338
rect 1582 2332 1585 2338
rect 1590 2302 1593 2348
rect 1630 2342 1633 2348
rect 1638 2332 1641 2418
rect 1670 2362 1673 2458
rect 1678 2452 1681 2498
rect 1726 2482 1729 2488
rect 1734 2482 1737 2528
rect 1750 2482 1753 2488
rect 1758 2482 1761 2528
rect 1782 2522 1785 2648
rect 1798 2592 1801 2658
rect 1806 2592 1809 2648
rect 1814 2632 1817 2668
rect 1822 2652 1825 2658
rect 1862 2652 1865 2698
rect 1834 2648 1838 2651
rect 1810 2568 1814 2571
rect 1790 2562 1793 2568
rect 1834 2558 1838 2561
rect 1862 2552 1865 2608
rect 1802 2548 1806 2551
rect 1818 2548 1822 2551
rect 1766 2492 1769 2498
rect 1790 2482 1793 2508
rect 1686 2472 1689 2478
rect 1694 2462 1697 2478
rect 1722 2468 1726 2471
rect 1710 2452 1713 2458
rect 1698 2438 1702 2441
rect 1742 2392 1745 2408
rect 1758 2392 1761 2468
rect 1730 2388 1734 2391
rect 1694 2352 1697 2358
rect 1658 2348 1662 2351
rect 1670 2342 1673 2348
rect 1718 2342 1721 2378
rect 1774 2362 1777 2468
rect 1790 2382 1793 2478
rect 1798 2462 1801 2538
rect 1838 2512 1841 2528
rect 1846 2522 1849 2528
rect 1814 2462 1817 2488
rect 1814 2411 1817 2458
rect 1810 2408 1817 2411
rect 1822 2432 1825 2448
rect 1822 2412 1825 2428
rect 1798 2362 1801 2398
rect 1818 2358 1822 2361
rect 1790 2352 1793 2358
rect 1830 2352 1833 2468
rect 1838 2462 1841 2508
rect 1862 2492 1865 2548
rect 1870 2491 1873 2868
rect 1918 2862 1921 3058
rect 1926 3052 1929 3138
rect 1942 3132 1945 3138
rect 1934 3082 1937 3108
rect 1934 3022 1937 3048
rect 1926 2952 1929 3018
rect 1942 2962 1945 3118
rect 1982 3102 1985 3118
rect 1990 3092 1993 3118
rect 1998 3082 2001 3158
rect 2014 3132 2017 3138
rect 2022 3122 2025 3158
rect 2042 3148 2046 3151
rect 2074 3148 2078 3151
rect 2046 3111 2049 3138
rect 2054 3122 2057 3138
rect 2066 3118 2070 3121
rect 2046 3108 2057 3111
rect 2054 3092 2057 3108
rect 2102 3092 2105 3148
rect 2126 3142 2129 3268
rect 2142 3262 2145 3338
rect 2194 3328 2198 3331
rect 2218 3318 2222 3321
rect 2182 3282 2185 3288
rect 2198 3202 2201 3268
rect 2254 3262 2257 3348
rect 2294 3332 2297 3388
rect 2342 3360 2345 3379
rect 2358 3372 2361 3418
rect 2454 3412 2457 3468
rect 2384 3403 2386 3407
rect 2390 3403 2393 3407
rect 2397 3403 2400 3407
rect 2394 3358 2398 3361
rect 2486 3352 2489 3458
rect 2526 3452 2529 3478
rect 2534 3462 2537 3468
rect 2542 3462 2545 3468
rect 2566 3462 2569 3488
rect 2578 3468 2582 3471
rect 2554 3458 2558 3461
rect 2570 3458 2574 3461
rect 2546 3448 2550 3451
rect 2502 3422 2505 3448
rect 2598 3422 2601 3448
rect 2526 3382 2529 3418
rect 2362 3348 2366 3351
rect 2310 3332 2313 3338
rect 2382 3322 2385 3338
rect 2526 3332 2529 3378
rect 2590 3362 2593 3388
rect 2294 3272 2297 3278
rect 2318 3272 2321 3308
rect 2338 3278 2342 3281
rect 2354 3278 2361 3281
rect 2302 3262 2305 3268
rect 2346 3258 2350 3261
rect 2230 3231 2233 3250
rect 2270 3232 2273 3248
rect 2286 3242 2289 3248
rect 2294 3212 2297 3258
rect 2310 3252 2313 3258
rect 2174 3192 2177 3198
rect 2294 3192 2297 3198
rect 2214 3162 2217 3168
rect 2226 3158 2230 3161
rect 2158 3152 2161 3158
rect 2122 3138 2126 3141
rect 2110 3132 2113 3138
rect 2134 3131 2137 3138
rect 2130 3128 2137 3131
rect 2118 3112 2121 3118
rect 2014 3082 2017 3088
rect 2066 3078 2073 3081
rect 1978 3068 1982 3071
rect 2042 3068 2046 3071
rect 2070 3071 2073 3078
rect 2070 3068 2086 3071
rect 2002 3058 2006 3061
rect 1986 3048 1990 3051
rect 1958 2942 1961 2988
rect 1954 2938 1958 2941
rect 1902 2831 1905 2850
rect 1906 2758 1910 2761
rect 1914 2748 1921 2751
rect 1894 2742 1897 2748
rect 1882 2738 1886 2741
rect 1910 2732 1913 2748
rect 1880 2703 1882 2707
rect 1886 2703 1889 2707
rect 1893 2703 1896 2707
rect 1902 2672 1905 2708
rect 1878 2662 1881 2668
rect 1890 2558 1894 2561
rect 1910 2552 1913 2718
rect 1918 2702 1921 2748
rect 1926 2672 1929 2858
rect 1942 2842 1945 2918
rect 1966 2892 1969 3048
rect 2014 2972 2017 3068
rect 2026 3058 2030 3061
rect 2038 3052 2041 3058
rect 2062 3052 2065 3068
rect 2118 3062 2121 3098
rect 2074 3058 2078 3061
rect 2126 3052 2129 3128
rect 2142 3072 2145 3148
rect 2170 3138 2174 3141
rect 2150 3062 2153 3098
rect 2190 3092 2193 3158
rect 2198 3152 2201 3158
rect 2218 3148 2222 3151
rect 2214 3092 2217 3138
rect 2222 3132 2225 3138
rect 2246 3132 2249 3138
rect 2234 3118 2238 3121
rect 2210 3078 2238 3081
rect 2174 3068 2182 3071
rect 2166 3062 2169 3068
rect 2138 3058 2142 3061
rect 2174 3061 2177 3068
rect 2170 3058 2177 3061
rect 2182 3052 2185 3058
rect 2198 3052 2201 3078
rect 2218 3068 2222 3071
rect 2246 3061 2249 3108
rect 2254 3102 2257 3138
rect 2262 3072 2265 3108
rect 2270 3082 2273 3158
rect 2294 3152 2297 3168
rect 2310 3142 2313 3208
rect 2326 3172 2329 3248
rect 2298 3138 2302 3141
rect 2318 3132 2321 3138
rect 2310 3092 2313 3108
rect 2302 3082 2305 3088
rect 2318 3081 2321 3108
rect 2310 3078 2321 3081
rect 2326 3082 2329 3138
rect 2334 3092 2337 3188
rect 2358 3172 2361 3278
rect 2370 3268 2374 3271
rect 2390 3262 2393 3318
rect 2402 3278 2406 3281
rect 2414 3272 2417 3318
rect 2422 3262 2425 3318
rect 2438 3282 2441 3328
rect 2446 3312 2449 3318
rect 2542 3312 2545 3338
rect 2590 3332 2593 3348
rect 2606 3332 2609 3458
rect 2494 3292 2497 3308
rect 2622 3292 2625 3408
rect 2646 3402 2649 3468
rect 2662 3422 2665 3478
rect 2702 3462 2705 3538
rect 2766 3532 2769 3578
rect 2902 3562 2905 3588
rect 2858 3548 2862 3551
rect 2890 3548 2894 3551
rect 2806 3542 2809 3548
rect 2910 3542 2913 3558
rect 2942 3552 2945 3588
rect 3118 3582 3121 3588
rect 2830 3492 2833 3528
rect 2850 3518 2854 3521
rect 2862 3492 2865 3528
rect 2886 3482 2889 3538
rect 2904 3503 2906 3507
rect 2910 3503 2913 3507
rect 2917 3503 2920 3507
rect 2926 3492 2929 3548
rect 2950 3542 2953 3568
rect 2990 3560 2993 3579
rect 3198 3572 3201 3578
rect 3230 3562 3233 3568
rect 2974 3542 2977 3548
rect 3150 3542 3153 3548
rect 3158 3542 3161 3558
rect 3174 3542 3177 3558
rect 3182 3552 3185 3558
rect 3226 3548 3230 3551
rect 3022 3532 3025 3538
rect 3038 3522 3041 3528
rect 3150 3522 3153 3528
rect 2902 3482 2905 3488
rect 2794 3468 2798 3471
rect 2858 3468 2862 3471
rect 2758 3452 2761 3458
rect 2746 3428 2750 3431
rect 2646 3360 2649 3379
rect 2774 3372 2777 3418
rect 2782 3372 2785 3418
rect 2638 3292 2641 3348
rect 2678 3342 2681 3348
rect 2678 3292 2681 3328
rect 2694 3302 2697 3328
rect 2442 3278 2446 3281
rect 2506 3278 2510 3281
rect 2522 3278 2526 3281
rect 2570 3278 2574 3281
rect 2514 3268 2518 3271
rect 2734 3271 2737 3348
rect 2786 3338 2790 3341
rect 2798 3322 2801 3458
rect 2814 3442 2817 3448
rect 2830 3412 2833 3458
rect 2846 3442 2849 3458
rect 2862 3342 2865 3448
rect 2878 3442 2881 3468
rect 2886 3452 2889 3458
rect 2934 3452 2937 3468
rect 2870 3382 2873 3438
rect 2870 3352 2873 3378
rect 2886 3362 2889 3448
rect 2878 3352 2881 3358
rect 2922 3348 2926 3351
rect 2886 3342 2889 3348
rect 2906 3338 2910 3341
rect 2782 3282 2785 3288
rect 2854 3282 2857 3338
rect 2734 3268 2745 3271
rect 2446 3262 2449 3268
rect 2598 3262 2601 3268
rect 2482 3258 2486 3261
rect 2546 3258 2550 3261
rect 2570 3258 2574 3261
rect 2366 3252 2369 3258
rect 2346 3158 2350 3161
rect 2366 3142 2369 3248
rect 2390 3242 2393 3248
rect 2374 3191 2377 3238
rect 2384 3203 2386 3207
rect 2390 3203 2393 3207
rect 2397 3203 2400 3207
rect 2374 3188 2385 3191
rect 2382 3162 2385 3188
rect 2414 3172 2417 3258
rect 2394 3168 2398 3171
rect 2414 3162 2417 3168
rect 2386 3158 2393 3161
rect 2362 3128 2366 3131
rect 2350 3092 2353 3128
rect 2298 3068 2302 3071
rect 2270 3062 2273 3068
rect 2242 3058 2249 3061
rect 2258 3058 2262 3061
rect 2282 3058 2286 3061
rect 2090 3048 2094 3051
rect 2234 3048 2238 3051
rect 1974 2962 1977 2968
rect 2030 2952 2033 2968
rect 1974 2842 1977 2918
rect 1982 2872 1985 2948
rect 2022 2942 2025 2948
rect 2002 2938 2006 2941
rect 1982 2852 1985 2858
rect 1942 2822 1945 2838
rect 1934 2752 1937 2768
rect 1942 2742 1945 2748
rect 1942 2682 1945 2738
rect 1954 2728 1958 2731
rect 1974 2722 1977 2838
rect 1990 2812 1993 2938
rect 2002 2928 2006 2931
rect 2014 2872 2017 2938
rect 2022 2872 2025 2878
rect 2014 2862 2017 2868
rect 1986 2768 1990 2771
rect 1998 2761 2001 2818
rect 2006 2792 2009 2818
rect 2022 2762 2025 2868
rect 1998 2758 2006 2761
rect 1986 2748 1990 2751
rect 2014 2742 2017 2758
rect 2030 2752 2033 2928
rect 2038 2902 2041 3048
rect 2102 3032 2105 3048
rect 2134 3042 2137 3048
rect 2046 2962 2049 2968
rect 2054 2962 2057 2978
rect 2062 2951 2065 2998
rect 2058 2948 2065 2951
rect 2070 2952 2073 3018
rect 2070 2932 2073 2938
rect 2062 2912 2065 2918
rect 2078 2912 2081 3018
rect 2094 2972 2097 2978
rect 2110 2962 2113 2998
rect 2126 2992 2129 3028
rect 2198 2972 2201 2978
rect 2142 2962 2145 2968
rect 2214 2962 2217 2968
rect 2162 2958 2177 2961
rect 2174 2951 2177 2958
rect 2174 2948 2182 2951
rect 2126 2942 2129 2948
rect 2134 2932 2137 2938
rect 2158 2922 2161 2948
rect 2222 2942 2225 2948
rect 2194 2938 2198 2941
rect 2182 2922 2185 2928
rect 2222 2922 2225 2928
rect 2046 2892 2049 2908
rect 2158 2902 2161 2918
rect 2070 2872 2073 2898
rect 2118 2892 2121 2898
rect 2098 2878 2102 2881
rect 2130 2878 2137 2881
rect 2134 2872 2137 2878
rect 2230 2872 2233 3048
rect 2270 3042 2273 3048
rect 2270 3022 2273 3038
rect 2262 2962 2265 2968
rect 2270 2952 2273 2958
rect 2310 2952 2313 3078
rect 2318 2962 2321 3058
rect 2342 3032 2345 3078
rect 2374 3072 2377 3148
rect 2390 3092 2393 3158
rect 2398 3152 2401 3158
rect 2422 3152 2425 3258
rect 2470 3252 2473 3258
rect 2590 3252 2593 3258
rect 2626 3248 2630 3251
rect 2438 3232 2441 3248
rect 2494 3242 2497 3248
rect 2438 3152 2441 3178
rect 2454 3142 2457 3148
rect 2442 3138 2446 3141
rect 2398 3102 2401 3138
rect 2466 3128 2470 3131
rect 2422 3082 2425 3088
rect 2362 3058 2366 3061
rect 2326 2972 2329 3018
rect 2334 2992 2337 2998
rect 2350 2982 2353 3048
rect 2246 2942 2249 2948
rect 2238 2882 2241 2938
rect 2258 2918 2262 2921
rect 2106 2868 2110 2871
rect 2194 2868 2198 2871
rect 2126 2862 2129 2868
rect 2150 2862 2153 2868
rect 2066 2858 2070 2861
rect 2082 2858 2086 2861
rect 2098 2858 2102 2861
rect 2138 2858 2142 2861
rect 2038 2852 2041 2858
rect 2158 2852 2161 2868
rect 2170 2858 2174 2861
rect 2210 2858 2214 2861
rect 2078 2812 2081 2848
rect 2166 2822 2169 2848
rect 2198 2842 2201 2848
rect 2222 2812 2225 2868
rect 2230 2862 2233 2868
rect 2078 2792 2081 2808
rect 2058 2748 2062 2751
rect 2038 2732 2041 2738
rect 2046 2732 2049 2738
rect 2070 2722 2073 2738
rect 2022 2712 2025 2718
rect 2094 2682 2097 2738
rect 2102 2682 2105 2808
rect 2222 2762 2225 2788
rect 2238 2782 2241 2878
rect 2250 2858 2254 2861
rect 2258 2848 2262 2851
rect 2110 2692 2113 2698
rect 1942 2632 1945 2678
rect 1998 2672 2001 2678
rect 1958 2662 1961 2668
rect 1922 2618 1926 2621
rect 1918 2542 1921 2608
rect 1942 2592 1945 2608
rect 1958 2552 1961 2658
rect 2014 2632 2017 2668
rect 2090 2658 2094 2661
rect 2062 2622 2065 2648
rect 2070 2560 2073 2579
rect 2094 2552 2097 2608
rect 1978 2548 1982 2551
rect 2102 2542 2105 2678
rect 2118 2672 2121 2758
rect 2174 2742 2177 2748
rect 2134 2692 2137 2708
rect 2158 2682 2161 2728
rect 2206 2692 2209 2728
rect 2214 2712 2217 2748
rect 2254 2742 2257 2848
rect 2262 2762 2265 2768
rect 2270 2762 2273 2938
rect 2294 2932 2297 2938
rect 2302 2932 2305 2948
rect 2282 2918 2286 2921
rect 2294 2872 2297 2908
rect 2302 2872 2305 2878
rect 2318 2872 2321 2958
rect 2350 2952 2353 2958
rect 2338 2948 2342 2951
rect 2366 2941 2369 3038
rect 2374 2972 2377 3068
rect 2382 3032 2385 3078
rect 2398 3062 2401 3068
rect 2422 3062 2425 3078
rect 2462 3071 2465 3118
rect 2478 3092 2481 3238
rect 2502 3192 2505 3248
rect 2566 3232 2569 3248
rect 2570 3228 2577 3231
rect 2510 3162 2513 3228
rect 2574 3162 2577 3228
rect 2514 3148 2518 3151
rect 2486 3092 2489 3148
rect 2514 3128 2518 3131
rect 2462 3068 2470 3071
rect 2438 3062 2441 3068
rect 2458 3058 2462 3061
rect 2430 3052 2433 3058
rect 2384 3003 2386 3007
rect 2390 3003 2393 3007
rect 2397 3003 2400 3007
rect 2414 2992 2417 3028
rect 2378 2948 2382 2951
rect 2366 2938 2377 2941
rect 2350 2932 2353 2938
rect 2342 2892 2345 2908
rect 2366 2892 2369 2928
rect 2374 2912 2377 2938
rect 2382 2932 2385 2938
rect 2398 2932 2401 2958
rect 2338 2868 2342 2871
rect 2278 2852 2281 2858
rect 2278 2772 2281 2818
rect 2286 2792 2289 2868
rect 2314 2848 2318 2851
rect 2302 2792 2305 2848
rect 2302 2782 2305 2788
rect 2286 2752 2289 2768
rect 2266 2748 2270 2751
rect 2294 2742 2297 2748
rect 2310 2741 2313 2758
rect 2318 2752 2321 2768
rect 2310 2738 2321 2741
rect 2286 2732 2289 2738
rect 2246 2712 2249 2718
rect 2218 2678 2222 2681
rect 2238 2672 2241 2678
rect 2246 2672 2249 2708
rect 2254 2672 2257 2678
rect 2138 2668 2142 2671
rect 2170 2668 2174 2671
rect 2218 2668 2222 2671
rect 2146 2658 2150 2661
rect 2110 2562 2113 2648
rect 2118 2572 2121 2658
rect 2166 2652 2169 2668
rect 2190 2662 2193 2668
rect 2114 2558 2118 2561
rect 2134 2552 2137 2568
rect 2150 2562 2153 2618
rect 2166 2592 2169 2648
rect 2142 2552 2145 2558
rect 1906 2538 1910 2541
rect 2122 2538 2126 2541
rect 1880 2503 1882 2507
rect 1886 2503 1889 2507
rect 1893 2503 1896 2507
rect 1926 2502 1929 2518
rect 1870 2488 1878 2491
rect 1846 2472 1849 2478
rect 1854 2472 1857 2478
rect 1894 2472 1897 2478
rect 1958 2472 1961 2498
rect 1894 2462 1897 2468
rect 1938 2458 1942 2461
rect 1846 2452 1849 2458
rect 1854 2452 1857 2458
rect 1926 2452 1929 2458
rect 1950 2402 1953 2468
rect 1966 2462 1969 2488
rect 1930 2358 1937 2361
rect 1870 2352 1873 2358
rect 1778 2348 1782 2351
rect 1850 2348 1854 2351
rect 1882 2348 1886 2351
rect 1806 2342 1809 2348
rect 1690 2338 1694 2341
rect 1714 2338 1718 2341
rect 1778 2338 1782 2341
rect 1662 2332 1665 2338
rect 1614 2282 1617 2328
rect 1638 2301 1641 2318
rect 1630 2298 1641 2301
rect 1630 2272 1633 2298
rect 1702 2292 1705 2328
rect 1734 2312 1737 2328
rect 1750 2282 1753 2328
rect 1766 2292 1769 2328
rect 1738 2268 1745 2271
rect 1570 2258 1574 2261
rect 1554 2158 1558 2161
rect 1566 2152 1569 2178
rect 1606 2142 1609 2148
rect 1614 2142 1617 2218
rect 1622 2162 1625 2198
rect 1630 2152 1633 2248
rect 1662 2231 1665 2250
rect 1698 2248 1702 2251
rect 1730 2248 1734 2251
rect 1742 2212 1745 2268
rect 1750 2262 1753 2268
rect 1646 2162 1649 2168
rect 1734 2162 1737 2208
rect 1662 2142 1665 2158
rect 1670 2142 1673 2148
rect 1634 2138 1638 2141
rect 1650 2138 1654 2141
rect 1582 2132 1585 2138
rect 1550 2062 1553 2128
rect 1582 2112 1585 2128
rect 1550 1981 1553 2028
rect 1542 1978 1553 1981
rect 1450 1938 1454 1941
rect 1390 1892 1393 1898
rect 1334 1862 1337 1868
rect 1360 1803 1362 1807
rect 1366 1803 1369 1807
rect 1373 1803 1376 1807
rect 1274 1788 1278 1791
rect 1246 1762 1249 1778
rect 1406 1772 1409 1938
rect 1414 1882 1417 1918
rect 1422 1852 1425 1888
rect 1434 1858 1438 1861
rect 1438 1842 1441 1848
rect 1374 1752 1377 1758
rect 1238 1692 1241 1708
rect 1246 1692 1249 1698
rect 1254 1682 1257 1718
rect 1262 1702 1265 1738
rect 1358 1732 1361 1738
rect 1374 1732 1377 1738
rect 1318 1692 1321 1718
rect 1374 1682 1377 1718
rect 1358 1672 1361 1678
rect 1234 1668 1238 1671
rect 1314 1668 1318 1671
rect 1190 1588 1201 1591
rect 1206 1638 1214 1641
rect 1166 1562 1169 1568
rect 1190 1562 1193 1588
rect 1198 1542 1201 1578
rect 1206 1572 1209 1638
rect 1230 1612 1233 1658
rect 1262 1642 1265 1668
rect 1334 1662 1337 1668
rect 1230 1592 1233 1598
rect 1270 1592 1273 1658
rect 1286 1622 1289 1648
rect 1342 1642 1345 1668
rect 1370 1658 1374 1661
rect 1106 1538 1110 1541
rect 1030 1532 1033 1538
rect 1046 1472 1049 1478
rect 1054 1472 1057 1528
rect 1114 1518 1118 1521
rect 1070 1472 1073 1518
rect 1094 1491 1097 1518
rect 1090 1488 1097 1491
rect 1102 1492 1105 1518
rect 1142 1512 1145 1518
rect 1150 1502 1153 1538
rect 1146 1488 1150 1491
rect 1166 1491 1169 1528
rect 1182 1512 1185 1528
rect 1166 1488 1174 1491
rect 1078 1478 1094 1481
rect 1154 1478 1161 1481
rect 998 1462 1001 1468
rect 950 1442 953 1448
rect 958 1432 961 1438
rect 946 1358 950 1361
rect 914 1348 918 1351
rect 930 1338 934 1341
rect 818 1258 822 1261
rect 830 1162 833 1328
rect 848 1303 850 1307
rect 854 1303 857 1307
rect 861 1303 864 1307
rect 870 1272 873 1318
rect 902 1312 905 1338
rect 918 1322 921 1338
rect 918 1312 921 1318
rect 926 1282 929 1318
rect 838 1231 841 1250
rect 886 1192 889 1278
rect 934 1222 937 1318
rect 846 1172 849 1178
rect 806 1142 809 1148
rect 614 1082 617 1088
rect 710 1082 713 1118
rect 782 1102 785 1138
rect 798 1112 801 1138
rect 830 1132 833 1158
rect 878 1152 881 1158
rect 842 1148 846 1151
rect 866 1148 870 1151
rect 822 1102 825 1118
rect 848 1103 850 1107
rect 854 1103 857 1107
rect 861 1103 864 1107
rect 742 1092 745 1098
rect 822 1082 825 1088
rect 566 1068 577 1071
rect 698 1068 702 1071
rect 398 872 401 888
rect 414 882 417 888
rect 446 872 449 878
rect 430 862 433 868
rect 454 862 457 888
rect 462 882 465 898
rect 470 882 473 938
rect 478 862 481 868
rect 486 862 489 938
rect 494 892 497 938
rect 502 862 505 898
rect 510 872 513 928
rect 526 902 529 938
rect 534 922 537 928
rect 530 888 534 891
rect 542 882 545 958
rect 566 942 569 1068
rect 574 1031 577 1058
rect 630 1032 633 1068
rect 710 1062 713 1078
rect 822 1072 825 1078
rect 838 1072 841 1098
rect 886 1072 889 1188
rect 894 1152 897 1198
rect 914 1168 918 1171
rect 902 1142 905 1158
rect 910 1142 913 1148
rect 926 1142 929 1148
rect 942 1142 945 1358
rect 958 1352 961 1418
rect 966 1352 969 1458
rect 978 1348 982 1351
rect 994 1348 998 1351
rect 1006 1342 1009 1468
rect 1030 1462 1033 1468
rect 1058 1458 1062 1461
rect 1078 1452 1081 1478
rect 1090 1468 1094 1471
rect 1138 1468 1142 1471
rect 1158 1471 1161 1478
rect 1190 1472 1193 1488
rect 1206 1472 1209 1548
rect 1158 1468 1174 1471
rect 954 1338 958 1341
rect 986 1338 990 1341
rect 950 1272 953 1338
rect 966 1292 969 1308
rect 974 1262 977 1318
rect 990 1292 993 1298
rect 998 1282 1001 1328
rect 1006 1292 1009 1318
rect 962 1148 966 1151
rect 898 1138 902 1141
rect 942 1122 945 1128
rect 942 1071 945 1118
rect 974 1092 977 1118
rect 982 1092 985 1278
rect 1022 1262 1025 1368
rect 1030 1302 1033 1438
rect 1086 1422 1089 1458
rect 1118 1402 1121 1458
rect 1038 1360 1041 1379
rect 1126 1372 1129 1458
rect 1130 1348 1134 1351
rect 1070 1342 1073 1348
rect 1086 1322 1089 1328
rect 1062 1308 1070 1311
rect 1062 1292 1065 1308
rect 1030 1272 1033 1288
rect 1086 1282 1089 1308
rect 1142 1302 1145 1468
rect 1150 1462 1153 1468
rect 1198 1462 1201 1468
rect 1222 1462 1225 1578
rect 1234 1468 1238 1471
rect 1166 1422 1169 1458
rect 1182 1452 1185 1458
rect 1166 1392 1169 1398
rect 1166 1372 1169 1388
rect 1198 1362 1201 1388
rect 1206 1352 1209 1448
rect 1222 1402 1225 1458
rect 1270 1452 1273 1548
rect 1310 1532 1313 1638
rect 1350 1612 1353 1658
rect 1360 1603 1362 1607
rect 1366 1603 1369 1607
rect 1373 1603 1376 1607
rect 1374 1562 1377 1588
rect 1326 1542 1329 1548
rect 1382 1542 1385 1658
rect 1398 1652 1401 1698
rect 1414 1672 1417 1768
rect 1422 1762 1425 1788
rect 1446 1762 1449 1818
rect 1454 1782 1457 1938
rect 1462 1932 1465 1958
rect 1494 1952 1497 1968
rect 1518 1952 1521 1958
rect 1474 1948 1478 1951
rect 1530 1928 1534 1931
rect 1486 1872 1489 1888
rect 1502 1871 1505 1918
rect 1510 1882 1513 1928
rect 1526 1892 1529 1918
rect 1534 1892 1537 1898
rect 1542 1872 1545 1978
rect 1558 1942 1561 2108
rect 1638 2072 1641 2078
rect 1582 2062 1585 2068
rect 1566 1992 1569 2038
rect 1590 2031 1593 2050
rect 1622 2042 1625 2068
rect 1694 2062 1697 2138
rect 1702 2132 1705 2158
rect 1726 2112 1729 2138
rect 1714 2088 1718 2091
rect 1718 2082 1721 2088
rect 1582 1962 1585 1968
rect 1590 1952 1593 1998
rect 1630 1972 1633 1978
rect 1654 1962 1657 2008
rect 1726 1992 1729 2068
rect 1742 2062 1745 2068
rect 1742 2042 1745 2048
rect 1750 2032 1753 2258
rect 1758 2252 1761 2288
rect 1782 2272 1785 2338
rect 1814 2332 1817 2348
rect 1838 2321 1841 2348
rect 1850 2338 1854 2341
rect 1850 2328 1854 2331
rect 1862 2328 1870 2331
rect 1838 2318 1849 2321
rect 1846 2292 1849 2318
rect 1862 2312 1865 2328
rect 1918 2322 1921 2348
rect 1870 2282 1873 2318
rect 1880 2303 1882 2307
rect 1886 2303 1889 2307
rect 1893 2303 1896 2307
rect 1862 2272 1865 2278
rect 1902 2272 1905 2318
rect 1934 2292 1937 2358
rect 1794 2268 1798 2271
rect 1818 2268 1822 2271
rect 1914 2268 1918 2271
rect 1774 2262 1777 2268
rect 1786 2248 1790 2251
rect 1774 2242 1777 2248
rect 1758 2152 1761 2238
rect 1814 2212 1817 2268
rect 1838 2262 1841 2268
rect 1826 2248 1838 2251
rect 1842 2248 1846 2251
rect 1862 2192 1865 2268
rect 1870 2262 1873 2268
rect 1766 2142 1769 2168
rect 1790 2152 1793 2178
rect 1818 2158 1822 2161
rect 1846 2152 1849 2158
rect 1802 2148 1806 2151
rect 1774 2142 1777 2148
rect 1766 2092 1769 2138
rect 1774 2102 1777 2138
rect 1766 2072 1769 2078
rect 1798 2072 1801 2138
rect 1806 2082 1809 2148
rect 1834 2138 1838 2141
rect 1862 2132 1865 2158
rect 1878 2142 1881 2258
rect 1878 2122 1881 2138
rect 1886 2132 1889 2258
rect 1926 2252 1929 2278
rect 1942 2272 1945 2348
rect 1974 2342 1977 2538
rect 1982 2452 1985 2518
rect 2014 2492 2017 2508
rect 2006 2472 2009 2478
rect 1994 2388 1998 2391
rect 1954 2338 1958 2341
rect 1974 2312 1977 2338
rect 1982 2332 1985 2358
rect 2006 2342 2009 2468
rect 2022 2422 2025 2528
rect 2038 2512 2041 2538
rect 2146 2528 2150 2531
rect 2054 2492 2057 2508
rect 2030 2462 2033 2478
rect 2038 2452 2041 2468
rect 2062 2462 2065 2478
rect 2074 2468 2078 2471
rect 2082 2458 2086 2461
rect 2046 2392 2049 2458
rect 2078 2442 2081 2448
rect 2026 2358 2030 2361
rect 2038 2352 2041 2388
rect 2026 2348 2030 2351
rect 2014 2342 2017 2348
rect 1986 2328 1990 2331
rect 1982 2292 1985 2318
rect 1998 2292 2001 2328
rect 1950 2262 1953 2268
rect 1902 2152 1905 2248
rect 1958 2222 1961 2268
rect 1974 2222 1977 2278
rect 1966 2192 1969 2218
rect 1918 2162 1921 2168
rect 1926 2151 1929 2188
rect 1950 2162 1953 2168
rect 1922 2148 1929 2151
rect 1962 2158 1966 2161
rect 1978 2158 1982 2161
rect 1914 2138 1918 2141
rect 1846 2092 1849 2118
rect 1934 2111 1937 2158
rect 1990 2152 1993 2288
rect 2014 2272 2017 2338
rect 2038 2302 2041 2338
rect 2046 2332 2049 2388
rect 2074 2368 2078 2371
rect 2062 2302 2065 2358
rect 2094 2272 2097 2528
rect 2102 2472 2105 2498
rect 2118 2462 2121 2518
rect 2158 2472 2161 2498
rect 2146 2468 2150 2471
rect 2118 2452 2121 2458
rect 2126 2442 2129 2458
rect 1998 2252 2001 2258
rect 2006 2232 2009 2248
rect 2022 2242 2025 2258
rect 2030 2252 2033 2268
rect 2094 2262 2097 2268
rect 2102 2262 2105 2438
rect 2158 2342 2161 2468
rect 2166 2462 2169 2548
rect 2182 2542 2185 2618
rect 2182 2492 2185 2518
rect 2190 2512 2193 2658
rect 2198 2472 2201 2668
rect 2230 2662 2233 2668
rect 2246 2652 2249 2658
rect 2262 2652 2265 2658
rect 2278 2622 2281 2648
rect 2310 2632 2313 2668
rect 2318 2662 2321 2738
rect 2318 2652 2321 2658
rect 2298 2628 2302 2631
rect 2206 2552 2209 2608
rect 2318 2592 2321 2648
rect 2262 2542 2265 2578
rect 2302 2532 2305 2588
rect 2310 2562 2313 2588
rect 2326 2552 2329 2858
rect 2334 2848 2342 2851
rect 2334 2762 2337 2848
rect 2342 2812 2345 2838
rect 2342 2762 2345 2808
rect 2366 2762 2369 2868
rect 2374 2852 2377 2908
rect 2398 2872 2401 2878
rect 2406 2872 2409 2968
rect 2430 2962 2433 2968
rect 2422 2942 2425 2948
rect 2430 2942 2433 2948
rect 2422 2882 2425 2888
rect 2386 2858 2390 2861
rect 2384 2803 2386 2807
rect 2390 2803 2393 2807
rect 2397 2803 2400 2807
rect 2370 2758 2374 2761
rect 2362 2748 2366 2751
rect 2342 2741 2345 2748
rect 2338 2738 2345 2741
rect 2342 2672 2345 2738
rect 2378 2738 2382 2741
rect 2366 2712 2369 2738
rect 2342 2641 2345 2668
rect 2350 2652 2353 2678
rect 2390 2672 2393 2788
rect 2414 2752 2417 2878
rect 2422 2792 2425 2868
rect 2438 2862 2441 3058
rect 2446 3042 2449 3048
rect 2462 3042 2465 3048
rect 2462 2992 2465 3008
rect 2462 2962 2465 2978
rect 2470 2962 2473 3068
rect 2478 3042 2481 3048
rect 2486 3022 2489 3088
rect 2494 3072 2497 3078
rect 2502 2982 2505 3068
rect 2510 3012 2513 3058
rect 2526 3052 2529 3158
rect 2566 3152 2569 3158
rect 2546 3148 2550 3151
rect 2578 3148 2582 3151
rect 2534 3102 2537 3148
rect 2566 3132 2569 3138
rect 2590 3102 2593 3248
rect 2646 3192 2649 3268
rect 2742 3262 2745 3268
rect 2798 3262 2801 3268
rect 2606 3162 2609 3168
rect 2622 3152 2625 3178
rect 2642 3148 2646 3151
rect 2602 3138 2606 3141
rect 2598 3092 2601 3118
rect 2630 3102 2633 3138
rect 2526 2972 2529 3048
rect 2534 3032 2537 3068
rect 2566 3062 2569 3078
rect 2622 3072 2625 3098
rect 2638 3091 2641 3138
rect 2634 3088 2641 3091
rect 2654 3082 2657 3258
rect 2674 3158 2681 3161
rect 2578 3068 2582 3071
rect 2590 3062 2593 3068
rect 2610 3058 2614 3061
rect 2566 3052 2569 3058
rect 2542 3032 2545 3038
rect 2566 2982 2569 3038
rect 2478 2962 2481 2968
rect 2542 2962 2545 2968
rect 2450 2958 2454 2961
rect 2450 2948 2454 2951
rect 2454 2892 2457 2938
rect 2462 2892 2465 2958
rect 2514 2948 2518 2951
rect 2478 2872 2481 2948
rect 2498 2938 2502 2941
rect 2534 2922 2537 2938
rect 2486 2892 2489 2918
rect 2542 2882 2545 2898
rect 2558 2872 2561 2948
rect 2566 2942 2569 2978
rect 2578 2938 2581 2941
rect 2582 2872 2585 2938
rect 2606 2912 2609 3048
rect 2622 2982 2625 3068
rect 2662 3062 2665 3098
rect 2670 3072 2673 3078
rect 2678 3072 2681 3158
rect 2686 3112 2689 3138
rect 2694 3092 2697 3248
rect 2702 3112 2705 3218
rect 2742 3202 2745 3258
rect 2830 3222 2833 3250
rect 2726 3160 2729 3179
rect 2758 3152 2761 3198
rect 2702 3072 2705 3108
rect 2666 3058 2670 3061
rect 2678 3052 2681 3068
rect 2710 3062 2713 3148
rect 2758 3132 2761 3138
rect 2774 3132 2777 3138
rect 2854 3082 2857 3278
rect 2862 3172 2865 3338
rect 2894 3332 2897 3338
rect 2870 3272 2873 3308
rect 2904 3303 2906 3307
rect 2910 3303 2913 3307
rect 2917 3303 2920 3307
rect 2898 3288 2902 3291
rect 2918 3272 2921 3278
rect 2926 3272 2929 3348
rect 2934 3332 2937 3418
rect 2950 3402 2953 3468
rect 2998 3462 3001 3498
rect 3014 3462 3017 3468
rect 3006 3452 3009 3458
rect 3014 3452 3017 3458
rect 3038 3452 3041 3488
rect 3078 3482 3081 3508
rect 3118 3492 3121 3518
rect 3150 3482 3153 3518
rect 3158 3512 3161 3538
rect 3158 3482 3161 3498
rect 3118 3472 3121 3478
rect 3054 3468 3062 3471
rect 2962 3448 2966 3451
rect 2982 3442 2985 3448
rect 2942 3398 2950 3401
rect 2942 3342 2945 3398
rect 2954 3388 2958 3391
rect 2950 3352 2953 3378
rect 2966 3362 2969 3418
rect 2966 3342 2969 3348
rect 2974 3332 2977 3438
rect 2982 3332 2985 3388
rect 2918 3152 2921 3248
rect 2926 3162 2929 3168
rect 2934 3152 2937 3328
rect 2950 3292 2953 3308
rect 2974 3292 2977 3328
rect 2982 3312 2985 3328
rect 2990 3282 2993 3408
rect 3022 3382 3025 3418
rect 3006 3362 3009 3378
rect 2998 3352 3001 3358
rect 3018 3348 3022 3351
rect 3030 3342 3033 3438
rect 2998 3332 3001 3338
rect 3014 3292 3017 3298
rect 3010 3278 3014 3281
rect 2954 3268 2958 3271
rect 2970 3268 2974 3271
rect 2958 3262 2961 3268
rect 2986 3258 2990 3261
rect 3014 3252 3017 3268
rect 3030 3262 3033 3308
rect 3038 3302 3041 3448
rect 3054 3362 3057 3468
rect 3074 3458 3078 3461
rect 3114 3458 3118 3461
rect 3062 3422 3065 3458
rect 3130 3448 3134 3451
rect 3142 3442 3145 3468
rect 3190 3462 3193 3508
rect 3174 3422 3177 3458
rect 3098 3368 3102 3371
rect 3110 3342 3113 3348
rect 3062 3322 3065 3332
rect 3038 3282 3041 3298
rect 3046 3272 3049 3318
rect 3022 3161 3025 3258
rect 3038 3242 3041 3268
rect 3054 3262 3057 3318
rect 3086 3312 3089 3338
rect 3098 3318 3102 3321
rect 3062 3252 3065 3258
rect 3054 3192 3057 3218
rect 3018 3158 3025 3161
rect 2998 3142 3001 3148
rect 3014 3142 3017 3148
rect 3022 3142 3025 3158
rect 3070 3152 3073 3298
rect 3078 3162 3081 3218
rect 3078 3142 3081 3158
rect 3086 3142 3089 3268
rect 3094 3252 3097 3278
rect 3110 3262 3113 3338
rect 3118 3292 3121 3358
rect 3126 3352 3129 3358
rect 3166 3352 3169 3418
rect 3190 3382 3193 3418
rect 3198 3392 3201 3548
rect 3210 3538 3214 3541
rect 3214 3452 3217 3488
rect 3230 3452 3233 3458
rect 3210 3448 3214 3451
rect 3222 3412 3225 3448
rect 3238 3442 3241 3578
rect 3262 3552 3265 3588
rect 3342 3582 3345 3588
rect 3482 3568 3486 3571
rect 3674 3568 3678 3571
rect 3318 3562 3321 3568
rect 3278 3552 3281 3558
rect 3246 3542 3249 3548
rect 3254 3532 3257 3538
rect 3254 3442 3257 3458
rect 3262 3442 3265 3508
rect 3278 3502 3281 3548
rect 3286 3542 3289 3548
rect 3326 3542 3329 3548
rect 3314 3538 3318 3541
rect 3294 3522 3297 3538
rect 3302 3528 3310 3531
rect 3294 3462 3297 3508
rect 3302 3482 3305 3528
rect 3334 3522 3337 3558
rect 3342 3511 3345 3568
rect 3390 3552 3393 3558
rect 3354 3548 3358 3551
rect 3426 3548 3430 3551
rect 3334 3508 3345 3511
rect 3334 3501 3337 3508
rect 3326 3498 3337 3501
rect 3310 3472 3313 3498
rect 3326 3471 3329 3498
rect 3318 3468 3329 3471
rect 3318 3461 3321 3468
rect 3350 3462 3353 3518
rect 3314 3458 3321 3461
rect 3330 3458 3337 3461
rect 3282 3448 3286 3451
rect 3234 3438 3238 3441
rect 3270 3422 3273 3448
rect 3242 3418 3246 3421
rect 3258 3418 3262 3421
rect 3222 3372 3225 3408
rect 3246 3392 3249 3418
rect 3258 3368 3262 3371
rect 3166 3342 3169 3348
rect 3138 3338 3142 3341
rect 3150 3292 3153 3328
rect 3118 3272 3121 3288
rect 3166 3282 3169 3338
rect 3174 3312 3177 3348
rect 3190 3342 3193 3368
rect 3206 3362 3209 3368
rect 3214 3352 3217 3368
rect 3222 3362 3225 3368
rect 3246 3362 3249 3368
rect 3278 3362 3281 3378
rect 3206 3322 3209 3328
rect 3174 3271 3177 3308
rect 3182 3282 3185 3318
rect 3174 3268 3182 3271
rect 3214 3271 3217 3348
rect 3230 3342 3233 3358
rect 3246 3342 3249 3358
rect 3270 3352 3273 3358
rect 3278 3352 3281 3358
rect 3230 3292 3233 3338
rect 3246 3302 3249 3338
rect 3270 3332 3273 3338
rect 3278 3312 3281 3348
rect 3246 3282 3249 3288
rect 3214 3268 3222 3271
rect 3126 3262 3129 3268
rect 3158 3262 3161 3268
rect 3114 3258 3121 3261
rect 3102 3252 3105 3258
rect 2862 3092 2865 3128
rect 2934 3122 2937 3138
rect 2990 3122 2993 3138
rect 3098 3128 3102 3131
rect 3110 3122 3113 3158
rect 2806 3072 2809 3078
rect 2698 3058 2702 3061
rect 2762 3058 2766 3061
rect 2646 3042 2649 3048
rect 2694 3042 2697 3048
rect 2710 2952 2713 3058
rect 2718 2982 2721 3038
rect 2822 3032 2825 3068
rect 2854 3022 2857 3050
rect 2726 3002 2729 3018
rect 2726 2962 2729 2988
rect 2622 2932 2625 2948
rect 2678 2942 2681 2948
rect 2750 2942 2753 2998
rect 2870 2952 2873 3058
rect 2878 3052 2881 3118
rect 2904 3103 2906 3107
rect 2910 3103 2913 3107
rect 2917 3103 2920 3107
rect 2974 3072 2977 3078
rect 2878 3022 2881 3048
rect 2902 2960 2905 2979
rect 2770 2938 2773 2941
rect 2662 2932 2665 2938
rect 2614 2892 2617 2918
rect 2662 2892 2665 2908
rect 2626 2878 2630 2881
rect 2646 2872 2649 2878
rect 2686 2872 2689 2908
rect 2742 2882 2745 2938
rect 2758 2892 2761 2918
rect 2766 2892 2769 2928
rect 2694 2872 2697 2878
rect 2774 2872 2777 2938
rect 2854 2932 2857 2938
rect 2870 2922 2873 2938
rect 2918 2922 2921 3018
rect 2926 2952 2929 2958
rect 2798 2892 2801 2908
rect 2904 2903 2906 2907
rect 2910 2903 2913 2907
rect 2917 2903 2920 2907
rect 2902 2882 2905 2888
rect 2810 2878 2814 2881
rect 2826 2878 2830 2881
rect 2610 2868 2614 2871
rect 2762 2868 2766 2871
rect 2438 2812 2441 2858
rect 2446 2822 2449 2858
rect 2462 2792 2465 2828
rect 2478 2792 2481 2868
rect 2570 2858 2574 2861
rect 2518 2852 2521 2858
rect 2590 2852 2593 2858
rect 2598 2852 2601 2858
rect 2622 2852 2625 2868
rect 2634 2858 2638 2861
rect 2662 2852 2665 2858
rect 2546 2848 2550 2851
rect 2650 2848 2654 2851
rect 2502 2842 2505 2848
rect 2518 2822 2521 2848
rect 2534 2812 2537 2818
rect 2590 2760 2593 2779
rect 2398 2732 2401 2738
rect 2414 2682 2417 2748
rect 2442 2738 2446 2741
rect 2422 2732 2425 2738
rect 2454 2732 2457 2748
rect 2438 2692 2441 2718
rect 2462 2692 2465 2698
rect 2446 2682 2449 2688
rect 2366 2662 2369 2668
rect 2342 2638 2361 2641
rect 2358 2562 2361 2638
rect 2374 2612 2377 2658
rect 2382 2652 2385 2668
rect 2418 2658 2422 2661
rect 2418 2648 2422 2651
rect 2430 2641 2433 2658
rect 2422 2638 2433 2641
rect 2446 2652 2449 2668
rect 2384 2603 2386 2607
rect 2390 2603 2393 2607
rect 2397 2603 2400 2607
rect 2406 2602 2409 2628
rect 2422 2592 2425 2638
rect 2386 2578 2390 2581
rect 2422 2572 2425 2588
rect 2446 2562 2449 2648
rect 2478 2562 2481 2758
rect 2542 2732 2545 2748
rect 2558 2732 2561 2738
rect 2598 2722 2601 2848
rect 2630 2762 2633 2768
rect 2606 2752 2609 2758
rect 2646 2752 2649 2818
rect 2678 2802 2681 2858
rect 2710 2852 2713 2858
rect 2690 2848 2694 2851
rect 2718 2842 2721 2868
rect 2662 2752 2665 2758
rect 2542 2672 2545 2678
rect 2370 2558 2374 2561
rect 2342 2542 2345 2548
rect 2334 2532 2337 2538
rect 2246 2522 2249 2528
rect 2230 2492 2233 2508
rect 2262 2492 2265 2528
rect 2282 2488 2286 2491
rect 2206 2482 2209 2488
rect 2222 2462 2225 2478
rect 2238 2462 2241 2488
rect 2310 2482 2313 2488
rect 2166 2392 2169 2458
rect 2182 2442 2185 2448
rect 2190 2432 2193 2458
rect 2222 2422 2225 2458
rect 2246 2432 2249 2458
rect 2286 2442 2289 2478
rect 2306 2468 2310 2471
rect 2318 2462 2321 2528
rect 2334 2492 2337 2518
rect 2350 2491 2353 2538
rect 2342 2488 2353 2491
rect 2342 2482 2345 2488
rect 2350 2462 2353 2478
rect 2262 2392 2265 2408
rect 2278 2402 2281 2418
rect 2358 2412 2361 2558
rect 2382 2552 2385 2558
rect 2426 2548 2430 2551
rect 2390 2522 2393 2538
rect 2406 2532 2409 2538
rect 2382 2492 2385 2508
rect 2406 2502 2409 2528
rect 2438 2522 2441 2558
rect 2454 2552 2457 2558
rect 2374 2482 2377 2488
rect 2422 2482 2425 2518
rect 2470 2502 2473 2538
rect 2366 2462 2369 2468
rect 2366 2442 2369 2448
rect 2222 2362 2225 2388
rect 2294 2382 2297 2388
rect 2306 2358 2310 2361
rect 2250 2348 2254 2351
rect 2282 2348 2286 2351
rect 2158 2322 2161 2328
rect 2174 2322 2177 2338
rect 2130 2268 2134 2271
rect 2170 2268 2174 2271
rect 2118 2262 2121 2268
rect 2222 2262 2225 2348
rect 2326 2342 2329 2348
rect 2314 2338 2318 2341
rect 2334 2332 2337 2338
rect 2366 2292 2369 2348
rect 2374 2292 2377 2478
rect 2390 2462 2393 2468
rect 2422 2452 2425 2478
rect 2430 2472 2433 2498
rect 2438 2468 2446 2471
rect 2438 2442 2441 2468
rect 2450 2458 2454 2461
rect 2470 2452 2473 2498
rect 2478 2452 2481 2558
rect 2494 2541 2497 2558
rect 2502 2552 2505 2638
rect 2558 2632 2561 2668
rect 2606 2662 2609 2748
rect 2694 2742 2697 2828
rect 2726 2772 2729 2858
rect 2734 2762 2737 2788
rect 2742 2752 2745 2758
rect 2714 2748 2718 2751
rect 2642 2738 2646 2741
rect 2666 2738 2670 2741
rect 2654 2722 2657 2738
rect 2686 2732 2689 2738
rect 2630 2672 2633 2698
rect 2638 2692 2641 2718
rect 2678 2702 2681 2718
rect 2646 2682 2649 2698
rect 2694 2681 2697 2738
rect 2702 2712 2705 2718
rect 2734 2692 2737 2728
rect 2694 2678 2702 2681
rect 2682 2668 2686 2671
rect 2694 2668 2702 2671
rect 2694 2662 2697 2668
rect 2590 2631 2593 2650
rect 2534 2592 2537 2598
rect 2510 2552 2513 2558
rect 2494 2538 2502 2541
rect 2514 2538 2518 2541
rect 2534 2532 2537 2558
rect 2542 2552 2545 2608
rect 2582 2572 2585 2578
rect 2598 2571 2601 2658
rect 2662 2652 2665 2658
rect 2718 2652 2721 2658
rect 2598 2568 2609 2571
rect 2550 2562 2553 2568
rect 2606 2562 2609 2568
rect 2638 2558 2646 2561
rect 2654 2561 2657 2648
rect 2742 2642 2745 2668
rect 2670 2632 2673 2638
rect 2750 2631 2753 2868
rect 2778 2858 2782 2861
rect 2774 2762 2777 2788
rect 2790 2772 2793 2818
rect 2814 2792 2817 2858
rect 2918 2812 2921 2868
rect 2950 2822 2953 2850
rect 2922 2788 2926 2791
rect 2794 2758 2801 2761
rect 2798 2752 2801 2758
rect 2786 2748 2790 2751
rect 2794 2738 2798 2741
rect 2766 2732 2769 2738
rect 2770 2728 2774 2731
rect 2758 2662 2761 2718
rect 2774 2662 2777 2698
rect 2794 2668 2798 2671
rect 2806 2671 2809 2738
rect 2822 2692 2825 2738
rect 2830 2732 2833 2758
rect 2862 2752 2865 2758
rect 2850 2748 2854 2751
rect 2874 2748 2878 2751
rect 2914 2748 2918 2751
rect 2850 2738 2854 2741
rect 2834 2728 2838 2731
rect 2802 2668 2809 2671
rect 2758 2642 2761 2648
rect 2742 2628 2753 2631
rect 2774 2632 2777 2638
rect 2670 2562 2673 2598
rect 2742 2592 2745 2628
rect 2782 2582 2785 2668
rect 2814 2662 2817 2668
rect 2798 2642 2801 2658
rect 2806 2592 2809 2628
rect 2814 2582 2817 2648
rect 2822 2642 2825 2648
rect 2830 2582 2833 2728
rect 2862 2702 2865 2748
rect 2850 2668 2854 2671
rect 2838 2592 2841 2658
rect 2702 2562 2705 2578
rect 2718 2562 2721 2568
rect 2654 2558 2662 2561
rect 2542 2522 2545 2538
rect 2534 2492 2537 2508
rect 2490 2478 2494 2481
rect 2384 2403 2386 2407
rect 2390 2403 2393 2407
rect 2397 2403 2400 2407
rect 2470 2402 2473 2448
rect 2390 2360 2393 2379
rect 2482 2348 2486 2351
rect 2422 2342 2425 2348
rect 2382 2292 2385 2338
rect 2438 2332 2441 2338
rect 2262 2282 2265 2288
rect 2046 2232 2049 2238
rect 2006 2212 2009 2228
rect 2014 2192 2017 2218
rect 2062 2201 2065 2258
rect 2102 2252 2105 2258
rect 2054 2198 2065 2201
rect 2158 2202 2161 2218
rect 1954 2148 1958 2151
rect 1970 2148 1974 2151
rect 1942 2112 1945 2138
rect 1934 2108 1942 2111
rect 1880 2103 1882 2107
rect 1886 2103 1889 2107
rect 1893 2103 1896 2107
rect 1870 2092 1873 2098
rect 1834 2078 1838 2081
rect 1866 2078 1870 2081
rect 1898 2078 1902 2081
rect 1966 2081 1969 2128
rect 1990 2102 1993 2148
rect 1998 2142 2001 2188
rect 2054 2182 2057 2198
rect 2222 2182 2225 2258
rect 2278 2221 2281 2268
rect 2326 2262 2329 2288
rect 2422 2282 2425 2328
rect 2494 2291 2497 2468
rect 2502 2442 2505 2458
rect 2510 2372 2513 2468
rect 2518 2382 2521 2418
rect 2534 2362 2537 2398
rect 2550 2362 2553 2508
rect 2566 2502 2569 2558
rect 2598 2552 2601 2558
rect 2638 2552 2641 2558
rect 2790 2552 2793 2558
rect 2578 2548 2582 2551
rect 2650 2548 2654 2551
rect 2666 2548 2670 2551
rect 2714 2548 2718 2551
rect 2746 2548 2753 2551
rect 2810 2548 2817 2551
rect 2574 2532 2577 2538
rect 2630 2522 2633 2538
rect 2638 2532 2641 2538
rect 2606 2502 2609 2518
rect 2614 2472 2617 2478
rect 2630 2472 2633 2498
rect 2686 2492 2689 2548
rect 2750 2542 2753 2548
rect 2738 2538 2742 2541
rect 2778 2538 2782 2541
rect 2802 2538 2806 2541
rect 2694 2472 2697 2538
rect 2726 2502 2729 2538
rect 2750 2492 2753 2538
rect 2766 2512 2769 2528
rect 2710 2472 2713 2478
rect 2754 2468 2758 2471
rect 2714 2458 2718 2461
rect 2550 2352 2553 2358
rect 2558 2342 2561 2378
rect 2538 2338 2542 2341
rect 2566 2332 2569 2368
rect 2574 2352 2577 2458
rect 2662 2431 2665 2450
rect 2586 2348 2590 2351
rect 2606 2342 2609 2358
rect 2518 2312 2521 2318
rect 2494 2288 2502 2291
rect 2358 2272 2361 2278
rect 2378 2268 2382 2271
rect 2414 2262 2417 2278
rect 2422 2272 2425 2278
rect 2462 2272 2465 2278
rect 2502 2272 2505 2288
rect 2514 2278 2518 2281
rect 2582 2272 2585 2298
rect 2590 2292 2593 2328
rect 2598 2322 2601 2328
rect 2614 2272 2617 2368
rect 2658 2358 2662 2361
rect 2634 2338 2638 2341
rect 2622 2272 2625 2328
rect 2646 2282 2649 2348
rect 2662 2342 2665 2348
rect 2654 2292 2657 2338
rect 2554 2268 2558 2271
rect 2446 2262 2449 2268
rect 2362 2258 2366 2261
rect 2310 2231 2313 2250
rect 2402 2248 2406 2251
rect 2278 2218 2289 2221
rect 2142 2160 2145 2179
rect 2158 2152 2161 2178
rect 2278 2162 2281 2168
rect 2230 2158 2238 2161
rect 2182 2152 2185 2158
rect 2202 2148 2206 2151
rect 2094 2132 2097 2138
rect 1974 2092 1977 2098
rect 1966 2078 1977 2081
rect 1786 2068 1790 2071
rect 1822 2052 1825 2058
rect 1762 2048 1766 2051
rect 1798 2048 1806 2051
rect 1782 2042 1785 2048
rect 1830 2042 1833 2068
rect 1774 2022 1777 2038
rect 1758 1972 1761 1978
rect 1710 1962 1713 1968
rect 1742 1962 1745 1968
rect 1774 1962 1777 2018
rect 1790 1992 1793 2028
rect 1606 1952 1609 1958
rect 1758 1952 1761 1958
rect 1666 1948 1670 1951
rect 1722 1948 1726 1951
rect 1566 1942 1569 1948
rect 1558 1932 1561 1938
rect 1550 1882 1553 1928
rect 1558 1892 1561 1908
rect 1574 1882 1577 1898
rect 1590 1892 1593 1938
rect 1502 1868 1510 1871
rect 1522 1868 1526 1871
rect 1586 1868 1590 1871
rect 1514 1858 1518 1861
rect 1478 1852 1481 1858
rect 1534 1842 1537 1848
rect 1526 1792 1529 1838
rect 1454 1742 1457 1768
rect 1478 1762 1481 1768
rect 1498 1758 1502 1761
rect 1542 1751 1545 1868
rect 1598 1861 1601 1948
rect 1630 1942 1633 1948
rect 1614 1932 1617 1938
rect 1622 1932 1625 1938
rect 1678 1902 1681 1938
rect 1686 1912 1689 1938
rect 1694 1922 1697 1948
rect 1782 1942 1785 1978
rect 1838 1972 1841 2078
rect 1874 2068 1878 2071
rect 1854 2032 1857 2058
rect 1862 1992 1865 2068
rect 1870 1982 1873 2068
rect 1886 2062 1889 2068
rect 1934 2062 1937 2068
rect 1942 2062 1945 2078
rect 1922 2058 1926 2061
rect 1906 2048 1910 2051
rect 1958 2032 1961 2058
rect 1810 1958 1814 1961
rect 1830 1952 1833 1958
rect 1818 1948 1822 1951
rect 1722 1938 1726 1941
rect 1718 1932 1721 1938
rect 1714 1918 1718 1921
rect 1646 1892 1649 1898
rect 1694 1892 1697 1908
rect 1750 1902 1753 1938
rect 1790 1912 1793 1948
rect 1822 1912 1825 1938
rect 1838 1932 1841 1968
rect 1846 1942 1849 1948
rect 1618 1888 1622 1891
rect 1790 1882 1793 1898
rect 1670 1872 1673 1878
rect 1806 1872 1809 1878
rect 1618 1868 1625 1871
rect 1598 1858 1606 1861
rect 1562 1838 1566 1841
rect 1550 1762 1553 1798
rect 1566 1762 1569 1768
rect 1574 1752 1577 1838
rect 1598 1832 1601 1848
rect 1598 1782 1601 1788
rect 1606 1782 1609 1858
rect 1582 1762 1585 1778
rect 1542 1748 1553 1751
rect 1414 1662 1417 1668
rect 1422 1592 1425 1688
rect 1454 1672 1457 1728
rect 1470 1702 1473 1718
rect 1486 1712 1489 1738
rect 1494 1722 1497 1738
rect 1506 1718 1510 1721
rect 1470 1678 1486 1681
rect 1462 1672 1465 1678
rect 1470 1672 1473 1678
rect 1430 1652 1433 1668
rect 1454 1582 1457 1668
rect 1462 1582 1465 1668
rect 1478 1652 1481 1668
rect 1494 1651 1497 1718
rect 1518 1711 1521 1738
rect 1526 1732 1529 1748
rect 1510 1708 1521 1711
rect 1502 1662 1505 1668
rect 1510 1661 1513 1708
rect 1518 1682 1521 1698
rect 1542 1692 1545 1728
rect 1526 1682 1529 1688
rect 1550 1672 1553 1748
rect 1594 1748 1598 1751
rect 1510 1658 1521 1661
rect 1490 1648 1497 1651
rect 1434 1568 1438 1571
rect 1470 1562 1473 1628
rect 1494 1592 1497 1638
rect 1518 1592 1521 1658
rect 1550 1612 1553 1668
rect 1522 1568 1526 1571
rect 1410 1558 1414 1561
rect 1506 1558 1510 1561
rect 1558 1552 1561 1748
rect 1606 1742 1609 1758
rect 1614 1752 1617 1848
rect 1622 1802 1625 1868
rect 1622 1752 1625 1758
rect 1570 1738 1574 1741
rect 1618 1738 1622 1741
rect 1606 1702 1609 1738
rect 1630 1712 1633 1868
rect 1638 1772 1641 1858
rect 1662 1852 1665 1858
rect 1646 1832 1649 1848
rect 1642 1758 1646 1761
rect 1642 1738 1646 1741
rect 1622 1672 1625 1698
rect 1638 1672 1641 1678
rect 1678 1672 1681 1868
rect 1854 1862 1857 1958
rect 1862 1922 1865 1938
rect 1862 1882 1865 1918
rect 1870 1892 1873 1948
rect 1926 1932 1929 2028
rect 1974 1992 1977 2078
rect 1990 1952 1993 1968
rect 2014 1962 2017 2058
rect 2026 1988 2030 1991
rect 2022 1952 2025 1958
rect 1962 1948 1966 1951
rect 1986 1938 1990 1941
rect 1914 1928 1918 1931
rect 1934 1912 1937 1938
rect 2030 1922 2033 1978
rect 2054 1942 2057 2078
rect 2070 2072 2073 2078
rect 2070 1952 2073 2058
rect 2102 2031 2105 2050
rect 2110 2042 2113 2138
rect 2150 2052 2153 2068
rect 2142 2012 2145 2018
rect 2158 1952 2161 2148
rect 2206 2132 2209 2138
rect 2190 2072 2193 2108
rect 2214 2082 2217 2158
rect 2230 2152 2233 2158
rect 2286 2151 2289 2218
rect 2298 2188 2302 2191
rect 2278 2148 2289 2151
rect 2294 2152 2297 2158
rect 2246 2142 2249 2148
rect 2222 2132 2225 2138
rect 2238 2092 2241 2138
rect 2226 2088 2230 2091
rect 2166 2062 2169 2068
rect 2222 2062 2225 2068
rect 2178 2048 2182 2051
rect 2174 1962 2177 1988
rect 2194 1958 2198 1961
rect 2206 1951 2209 2058
rect 2218 2048 2222 2051
rect 2230 1962 2233 2018
rect 2246 1992 2249 2138
rect 2254 2132 2257 2138
rect 2262 2062 2265 2118
rect 2270 2102 2273 2128
rect 2278 2092 2281 2148
rect 2310 2142 2313 2148
rect 2318 2142 2321 2188
rect 2302 2092 2305 2138
rect 2294 2082 2297 2088
rect 2326 2082 2329 2218
rect 2350 2212 2353 2248
rect 2342 2162 2345 2208
rect 2358 2152 2361 2248
rect 2384 2203 2386 2207
rect 2390 2203 2393 2207
rect 2397 2203 2400 2207
rect 2374 2172 2377 2198
rect 2430 2192 2433 2248
rect 2442 2238 2446 2241
rect 2454 2212 2457 2268
rect 2486 2262 2489 2268
rect 2494 2262 2497 2268
rect 2546 2258 2550 2261
rect 2578 2258 2582 2261
rect 2470 2242 2473 2258
rect 2590 2251 2593 2268
rect 2638 2262 2641 2268
rect 2610 2258 2614 2261
rect 2626 2258 2630 2261
rect 2582 2248 2593 2251
rect 2462 2182 2465 2188
rect 2486 2182 2489 2248
rect 2494 2192 2497 2238
rect 2374 2162 2377 2168
rect 2394 2158 2401 2161
rect 2398 2152 2401 2158
rect 2346 2148 2353 2151
rect 2342 2132 2345 2138
rect 2334 2102 2337 2128
rect 2350 2101 2353 2148
rect 2358 2142 2361 2148
rect 2390 2142 2393 2148
rect 2434 2138 2438 2141
rect 2366 2132 2369 2138
rect 2350 2098 2361 2101
rect 2358 2092 2361 2098
rect 2414 2092 2417 2138
rect 2422 2112 2425 2138
rect 2446 2132 2449 2158
rect 2462 2152 2465 2158
rect 2346 2088 2350 2091
rect 2306 2078 2310 2081
rect 2346 2078 2350 2081
rect 2270 1982 2273 2068
rect 2286 2062 2289 2078
rect 2302 2072 2305 2078
rect 2326 2072 2329 2078
rect 2306 2058 2310 2061
rect 2266 1958 2270 1961
rect 2278 1952 2281 2008
rect 2294 2002 2297 2018
rect 2326 2012 2329 2058
rect 2366 2031 2369 2058
rect 2390 2042 2393 2068
rect 2398 2062 2401 2088
rect 2378 2038 2382 2041
rect 2366 2028 2377 2031
rect 2374 2012 2377 2028
rect 2406 2012 2409 2078
rect 2454 2072 2457 2138
rect 2470 2132 2473 2178
rect 2478 2162 2481 2168
rect 2518 2162 2521 2188
rect 2506 2158 2510 2161
rect 2494 2152 2497 2158
rect 2482 2138 2486 2141
rect 2470 2092 2473 2128
rect 2518 2122 2521 2128
rect 2526 2112 2529 2248
rect 2558 2192 2561 2218
rect 2582 2192 2585 2248
rect 2622 2242 2625 2248
rect 2534 2152 2537 2158
rect 2554 2138 2561 2141
rect 2550 2122 2553 2128
rect 2502 2092 2505 2108
rect 2558 2092 2561 2138
rect 2566 2132 2569 2148
rect 2582 2092 2585 2118
rect 2606 2092 2609 2148
rect 2470 2072 2473 2088
rect 2326 1972 2329 1978
rect 2338 1958 2342 1961
rect 2350 1952 2353 1998
rect 2366 1952 2369 1958
rect 2206 1948 2214 1951
rect 2266 1948 2270 1951
rect 2126 1942 2129 1948
rect 2198 1942 2201 1948
rect 2110 1932 2113 1938
rect 2230 1932 2233 1948
rect 2246 1922 2249 1938
rect 2254 1932 2257 1948
rect 2286 1932 2289 1938
rect 1880 1903 1882 1907
rect 1886 1903 1889 1907
rect 1893 1903 1896 1907
rect 1950 1882 1953 1918
rect 1894 1872 1897 1878
rect 1930 1868 1934 1871
rect 1954 1868 1958 1871
rect 1694 1792 1697 1848
rect 1710 1822 1713 1848
rect 1838 1822 1841 1850
rect 1710 1802 1713 1818
rect 1694 1762 1697 1788
rect 1742 1752 1745 1778
rect 1782 1762 1785 1778
rect 1814 1762 1817 1818
rect 1750 1752 1753 1758
rect 1798 1752 1801 1758
rect 1830 1752 1833 1798
rect 1894 1762 1897 1828
rect 1902 1752 1905 1858
rect 1914 1848 1918 1851
rect 1918 1782 1921 1848
rect 1958 1842 1961 1848
rect 1930 1768 1934 1771
rect 1842 1748 1846 1751
rect 1726 1742 1729 1748
rect 1830 1742 1833 1748
rect 1570 1658 1574 1661
rect 1590 1631 1593 1650
rect 1574 1592 1577 1618
rect 1630 1592 1633 1598
rect 1598 1582 1601 1588
rect 1630 1552 1633 1588
rect 1710 1572 1713 1738
rect 1758 1732 1761 1738
rect 1750 1692 1753 1728
rect 1766 1692 1769 1718
rect 1774 1712 1777 1728
rect 1782 1722 1785 1728
rect 1806 1702 1809 1738
rect 1838 1732 1841 1738
rect 1814 1722 1817 1728
rect 1854 1722 1857 1738
rect 1910 1732 1913 1738
rect 1918 1732 1921 1738
rect 1926 1732 1929 1748
rect 1950 1732 1953 1748
rect 1790 1692 1793 1698
rect 1838 1692 1841 1698
rect 1818 1678 1822 1681
rect 1726 1672 1729 1678
rect 1778 1668 1782 1671
rect 1734 1592 1737 1668
rect 1758 1622 1761 1668
rect 1766 1662 1769 1668
rect 1846 1662 1849 1668
rect 1854 1662 1857 1678
rect 1778 1658 1782 1661
rect 1810 1658 1814 1661
rect 1458 1548 1462 1551
rect 1610 1548 1614 1551
rect 1430 1542 1433 1548
rect 1446 1532 1449 1538
rect 1494 1532 1497 1548
rect 1310 1511 1313 1528
rect 1310 1508 1321 1511
rect 1286 1492 1289 1508
rect 1302 1472 1305 1478
rect 1318 1472 1321 1508
rect 1326 1492 1329 1528
rect 1342 1482 1345 1508
rect 1502 1502 1505 1538
rect 1526 1512 1529 1548
rect 1558 1542 1561 1548
rect 1542 1522 1545 1528
rect 1362 1488 1366 1491
rect 1366 1472 1369 1488
rect 1310 1392 1313 1458
rect 1034 1258 1038 1261
rect 998 1252 1001 1258
rect 990 1152 993 1218
rect 1006 1192 1009 1248
rect 1022 1202 1025 1258
rect 1054 1192 1057 1278
rect 1102 1272 1105 1298
rect 1114 1268 1118 1271
rect 1126 1262 1129 1288
rect 1142 1282 1145 1288
rect 1154 1278 1158 1281
rect 1154 1268 1158 1271
rect 1178 1268 1182 1271
rect 1206 1262 1209 1348
rect 1246 1342 1249 1348
rect 1262 1322 1265 1328
rect 1254 1272 1257 1298
rect 1138 1258 1142 1261
rect 1086 1192 1089 1258
rect 1014 1152 1017 1158
rect 1054 1152 1057 1158
rect 1110 1152 1113 1228
rect 1074 1148 1078 1151
rect 1046 1142 1049 1148
rect 994 1138 998 1141
rect 1034 1138 1038 1141
rect 1082 1138 1086 1141
rect 1102 1132 1105 1138
rect 1106 1128 1113 1131
rect 1030 1122 1033 1128
rect 982 1081 985 1088
rect 978 1078 985 1081
rect 942 1068 953 1071
rect 722 1058 726 1061
rect 778 1058 782 1061
rect 938 1058 942 1061
rect 678 1042 681 1048
rect 574 992 577 998
rect 718 962 721 988
rect 750 952 753 1058
rect 950 1052 953 1068
rect 958 1062 961 1068
rect 974 1062 977 1078
rect 998 1072 1001 1078
rect 982 1062 985 1068
rect 990 1052 993 1068
rect 1006 1052 1009 1118
rect 1014 1062 1017 1068
rect 1022 1062 1025 1098
rect 1030 1072 1033 1078
rect 1030 1062 1033 1068
rect 870 1031 873 1050
rect 962 1048 966 1051
rect 902 992 905 1048
rect 930 1038 934 1041
rect 758 962 761 988
rect 926 962 929 1018
rect 998 1002 1001 1018
rect 950 952 953 998
rect 998 960 1001 979
rect 754 948 758 951
rect 914 948 918 951
rect 670 942 673 948
rect 550 892 553 918
rect 538 878 542 881
rect 394 858 398 861
rect 406 852 409 858
rect 378 838 382 841
rect 344 803 346 807
rect 350 803 353 807
rect 357 803 360 807
rect 390 792 393 818
rect 370 768 374 771
rect 406 752 409 848
rect 422 842 425 858
rect 338 728 342 731
rect 358 682 361 748
rect 386 728 390 731
rect 398 701 401 748
rect 406 712 409 748
rect 422 732 425 768
rect 470 761 473 818
rect 510 812 513 868
rect 494 792 497 808
rect 466 758 473 761
rect 486 752 489 758
rect 450 748 465 751
rect 462 742 465 748
rect 502 742 505 748
rect 482 738 486 741
rect 418 718 422 721
rect 398 698 406 701
rect 386 688 390 691
rect 326 672 329 678
rect 398 672 401 678
rect 394 658 398 661
rect 344 603 346 607
rect 350 603 353 607
rect 357 603 360 607
rect 374 592 377 658
rect 394 648 398 651
rect 406 641 409 698
rect 422 682 425 688
rect 398 638 409 641
rect 414 672 417 678
rect 430 671 433 718
rect 430 668 438 671
rect 398 592 401 638
rect 310 552 313 588
rect 402 568 406 571
rect 366 562 369 568
rect 390 542 393 558
rect 274 538 278 541
rect 362 538 366 541
rect 334 522 337 528
rect 382 502 385 538
rect 398 502 401 548
rect 414 532 417 668
rect 446 662 449 678
rect 454 672 457 738
rect 466 728 470 731
rect 422 562 425 658
rect 422 552 425 558
rect 430 542 433 618
rect 446 572 449 618
rect 366 492 369 498
rect 406 492 409 528
rect 422 522 425 538
rect 430 522 433 528
rect 294 472 297 478
rect 286 462 289 468
rect 258 458 262 461
rect 38 362 41 450
rect 126 431 129 458
rect 90 358 94 361
rect 38 254 41 358
rect 142 352 145 378
rect 70 302 73 338
rect 142 332 145 338
rect 86 282 89 298
rect 70 272 73 278
rect 86 192 89 278
rect 126 231 129 258
rect 110 192 113 208
rect 158 192 161 328
rect 170 288 174 291
rect 90 148 94 151
rect 6 142 9 148
rect 22 131 25 148
rect 34 138 38 141
rect 22 128 30 131
rect 118 92 121 188
rect 166 142 169 148
rect 118 82 121 88
rect 134 72 137 108
rect 6 42 9 48
rect 174 -19 177 118
rect 182 62 185 258
rect 190 152 193 218
rect 198 142 201 148
rect 222 62 225 218
rect 230 92 233 458
rect 266 448 270 451
rect 238 392 241 448
rect 262 392 265 438
rect 286 332 289 458
rect 294 452 297 458
rect 302 452 305 488
rect 394 468 398 471
rect 318 442 321 468
rect 326 462 329 468
rect 342 462 345 468
rect 414 462 417 468
rect 422 462 425 508
rect 438 462 441 568
rect 454 542 457 668
rect 462 652 465 708
rect 510 682 513 748
rect 486 672 489 678
rect 474 668 478 671
rect 474 658 478 661
rect 462 552 465 648
rect 510 592 513 678
rect 526 672 529 728
rect 550 692 553 868
rect 558 862 561 878
rect 558 742 561 818
rect 566 772 569 928
rect 654 922 657 928
rect 574 852 577 888
rect 590 882 593 888
rect 650 868 654 871
rect 702 862 705 948
rect 806 942 809 948
rect 1030 942 1033 948
rect 1046 942 1049 1018
rect 1086 952 1089 1098
rect 1094 1042 1097 1128
rect 1102 1072 1105 1078
rect 1110 1072 1113 1128
rect 1118 1071 1121 1258
rect 1134 1151 1137 1258
rect 1130 1148 1137 1151
rect 1158 1142 1161 1218
rect 1182 1202 1185 1258
rect 1166 1192 1169 1198
rect 1190 1162 1193 1168
rect 1158 1122 1161 1128
rect 1126 1082 1129 1118
rect 1166 1092 1169 1098
rect 1118 1068 1129 1071
rect 1102 962 1105 1068
rect 1114 1058 1118 1061
rect 1126 1052 1129 1068
rect 1142 1062 1145 1068
rect 1150 1062 1153 1078
rect 1190 1062 1193 1158
rect 1206 1152 1209 1258
rect 1270 1252 1273 1278
rect 1222 1231 1225 1250
rect 1294 1160 1297 1179
rect 1206 1102 1209 1148
rect 1246 1132 1249 1138
rect 1262 1122 1265 1138
rect 1318 1122 1321 1468
rect 1330 1458 1334 1461
rect 1350 1391 1353 1468
rect 1360 1403 1362 1407
rect 1366 1403 1369 1407
rect 1373 1403 1376 1407
rect 1350 1388 1358 1391
rect 1346 1328 1350 1331
rect 1370 1328 1374 1331
rect 1382 1292 1385 1388
rect 1390 1322 1393 1338
rect 1398 1292 1401 1498
rect 1446 1482 1449 1488
rect 1406 1452 1409 1458
rect 1462 1422 1465 1468
rect 1510 1422 1513 1448
rect 1446 1382 1449 1408
rect 1478 1382 1481 1388
rect 1446 1362 1449 1378
rect 1410 1358 1414 1361
rect 1438 1352 1441 1358
rect 1426 1348 1430 1351
rect 1406 1342 1409 1348
rect 1438 1332 1441 1338
rect 1446 1312 1449 1358
rect 1458 1348 1462 1351
rect 1486 1342 1489 1368
rect 1470 1302 1473 1318
rect 1446 1292 1449 1298
rect 1354 1278 1358 1281
rect 1390 1272 1393 1278
rect 1360 1203 1362 1207
rect 1366 1203 1369 1207
rect 1373 1203 1376 1207
rect 1390 1162 1393 1168
rect 1398 1151 1401 1288
rect 1470 1282 1473 1298
rect 1410 1278 1414 1281
rect 1454 1272 1457 1278
rect 1434 1258 1438 1261
rect 1406 1252 1409 1258
rect 1418 1158 1422 1161
rect 1446 1152 1449 1178
rect 1398 1148 1406 1151
rect 1470 1142 1473 1278
rect 1494 1262 1497 1358
rect 1502 1352 1505 1358
rect 1510 1352 1513 1368
rect 1526 1352 1529 1498
rect 1558 1472 1561 1538
rect 1710 1532 1713 1568
rect 1774 1562 1777 1588
rect 1766 1552 1769 1558
rect 1814 1552 1817 1658
rect 1726 1532 1729 1538
rect 1534 1462 1537 1468
rect 1554 1458 1557 1461
rect 1566 1452 1569 1528
rect 1582 1522 1585 1528
rect 1638 1452 1641 1478
rect 1654 1472 1657 1488
rect 1742 1472 1745 1498
rect 1766 1472 1769 1548
rect 1798 1532 1801 1548
rect 1786 1488 1790 1491
rect 1806 1472 1809 1488
rect 1822 1472 1825 1658
rect 1862 1651 1865 1718
rect 1870 1712 1873 1728
rect 1880 1703 1882 1707
rect 1886 1703 1889 1707
rect 1893 1703 1896 1707
rect 1870 1662 1873 1678
rect 1862 1648 1873 1651
rect 1870 1642 1873 1648
rect 1858 1638 1862 1641
rect 1834 1538 1838 1541
rect 1834 1528 1838 1531
rect 1834 1488 1838 1491
rect 1542 1362 1545 1418
rect 1566 1392 1569 1418
rect 1530 1348 1534 1351
rect 1518 1322 1521 1338
rect 1526 1332 1529 1338
rect 1550 1332 1553 1358
rect 1502 1262 1505 1268
rect 1494 1192 1497 1258
rect 1510 1251 1513 1308
rect 1534 1282 1537 1318
rect 1542 1292 1545 1328
rect 1506 1248 1513 1251
rect 1330 1138 1334 1141
rect 1354 1138 1358 1141
rect 1342 1132 1345 1138
rect 1222 1062 1225 1078
rect 1230 1072 1233 1078
rect 1238 1062 1241 1108
rect 1278 1092 1281 1108
rect 1262 1072 1265 1078
rect 1334 1072 1337 1118
rect 1342 1072 1345 1078
rect 1262 1062 1265 1068
rect 1126 992 1129 1048
rect 1134 1032 1137 1058
rect 1214 1052 1217 1058
rect 1254 1051 1257 1058
rect 1374 1052 1377 1058
rect 1382 1052 1385 1118
rect 1398 1062 1401 1138
rect 1414 1132 1417 1138
rect 1438 1132 1441 1138
rect 1478 1132 1481 1188
rect 1494 1152 1497 1188
rect 1462 1122 1465 1128
rect 1254 1048 1265 1051
rect 1354 1048 1358 1051
rect 954 938 958 941
rect 822 912 825 928
rect 1046 922 1049 928
rect 848 903 850 907
rect 854 903 857 907
rect 861 903 864 907
rect 930 888 934 891
rect 742 882 745 888
rect 1006 882 1009 888
rect 1022 872 1025 878
rect 850 868 854 871
rect 666 818 670 821
rect 638 752 641 778
rect 678 760 681 761
rect 674 756 678 759
rect 638 732 641 738
rect 622 722 625 728
rect 582 672 585 698
rect 606 692 609 708
rect 522 658 526 661
rect 510 562 513 568
rect 502 552 505 558
rect 522 548 526 551
rect 534 542 537 668
rect 586 658 590 661
rect 642 658 646 661
rect 546 588 550 591
rect 522 538 526 541
rect 478 482 481 528
rect 474 478 478 481
rect 446 472 449 478
rect 486 472 489 538
rect 494 492 497 518
rect 494 472 497 488
rect 514 468 518 471
rect 330 448 334 451
rect 382 442 385 458
rect 438 452 441 458
rect 398 442 401 448
rect 344 403 346 407
rect 350 403 353 407
rect 357 403 360 407
rect 446 391 449 468
rect 462 462 465 468
rect 542 462 545 548
rect 550 472 553 578
rect 558 572 561 648
rect 498 458 502 461
rect 454 452 457 458
rect 518 452 521 458
rect 542 452 545 458
rect 510 442 513 448
rect 526 442 529 448
rect 446 388 454 391
rect 310 362 313 368
rect 358 352 361 378
rect 486 362 489 388
rect 494 342 497 418
rect 358 332 361 338
rect 286 292 289 328
rect 270 212 273 278
rect 286 272 289 278
rect 338 258 342 261
rect 374 252 377 328
rect 502 312 505 348
rect 534 342 537 348
rect 550 342 553 468
rect 558 462 561 568
rect 590 552 593 658
rect 630 572 633 618
rect 646 552 649 578
rect 678 560 681 756
rect 702 712 705 858
rect 758 812 761 868
rect 790 831 793 850
rect 790 792 793 808
rect 902 792 905 868
rect 1086 862 1089 948
rect 1134 881 1137 1018
rect 1166 1012 1169 1018
rect 1198 962 1201 1018
rect 1206 992 1209 1048
rect 1238 992 1241 998
rect 1142 942 1145 948
rect 1150 942 1153 958
rect 1206 952 1209 988
rect 1162 948 1166 951
rect 1174 892 1177 948
rect 1182 932 1185 938
rect 1222 912 1225 928
rect 1134 878 1142 881
rect 1190 872 1193 908
rect 1198 882 1201 888
rect 1154 868 1158 871
rect 1210 868 1214 871
rect 1126 862 1129 868
rect 1134 862 1137 868
rect 1222 862 1225 888
rect 1254 882 1257 1018
rect 1262 982 1265 1048
rect 1278 952 1281 1008
rect 1360 1003 1362 1007
rect 1366 1003 1369 1007
rect 1373 1003 1376 1007
rect 1382 962 1385 988
rect 1390 952 1393 1058
rect 1398 1002 1401 1058
rect 1414 1052 1417 1058
rect 1430 1012 1433 1118
rect 1478 1112 1481 1128
rect 1494 1122 1497 1138
rect 1510 1082 1513 1238
rect 1518 1222 1521 1258
rect 1526 1252 1529 1268
rect 1534 1242 1537 1278
rect 1558 1271 1561 1348
rect 1566 1302 1569 1348
rect 1574 1342 1577 1368
rect 1598 1361 1601 1428
rect 1598 1358 1606 1361
rect 1594 1328 1598 1331
rect 1554 1268 1561 1271
rect 1566 1272 1569 1278
rect 1582 1262 1585 1278
rect 1614 1272 1617 1398
rect 1622 1332 1625 1348
rect 1630 1342 1633 1358
rect 1638 1352 1641 1418
rect 1646 1372 1649 1378
rect 1666 1358 1670 1361
rect 1686 1352 1689 1468
rect 1702 1462 1705 1468
rect 1726 1462 1729 1468
rect 1758 1462 1761 1468
rect 1774 1452 1777 1468
rect 1810 1458 1814 1461
rect 1702 1422 1705 1448
rect 1710 1382 1713 1388
rect 1718 1351 1721 1388
rect 1714 1348 1721 1351
rect 1638 1342 1641 1348
rect 1558 1252 1561 1258
rect 1518 1182 1521 1218
rect 1546 1168 1550 1171
rect 1570 1158 1574 1161
rect 1518 1142 1521 1158
rect 1546 1148 1550 1151
rect 1570 1148 1574 1151
rect 1534 1141 1537 1148
rect 1534 1138 1545 1141
rect 1530 1128 1534 1131
rect 1542 1122 1545 1138
rect 1558 1082 1561 1138
rect 1582 1121 1585 1258
rect 1598 1252 1601 1268
rect 1606 1262 1609 1268
rect 1598 1191 1601 1248
rect 1590 1188 1601 1191
rect 1590 1141 1593 1188
rect 1614 1171 1617 1268
rect 1638 1262 1641 1328
rect 1646 1292 1649 1348
rect 1686 1322 1689 1348
rect 1702 1342 1705 1348
rect 1694 1302 1697 1338
rect 1726 1312 1729 1348
rect 1734 1342 1737 1418
rect 1742 1372 1745 1378
rect 1750 1362 1753 1418
rect 1790 1392 1793 1458
rect 1798 1452 1801 1458
rect 1766 1362 1769 1378
rect 1774 1362 1777 1368
rect 1766 1352 1769 1358
rect 1786 1348 1790 1351
rect 1758 1342 1761 1348
rect 1798 1342 1801 1418
rect 1814 1411 1817 1448
rect 1822 1422 1825 1468
rect 1846 1452 1849 1578
rect 1878 1552 1881 1678
rect 1894 1662 1897 1688
rect 1902 1672 1905 1718
rect 1918 1682 1921 1688
rect 1926 1672 1929 1708
rect 1934 1692 1937 1698
rect 1942 1682 1945 1708
rect 1950 1682 1953 1728
rect 1914 1658 1918 1661
rect 1886 1652 1889 1658
rect 1886 1552 1889 1608
rect 1942 1592 1945 1678
rect 1958 1662 1961 1758
rect 1966 1742 1969 1878
rect 1974 1762 1977 1918
rect 2030 1872 2033 1918
rect 2038 1882 2041 1888
rect 2090 1878 2094 1881
rect 1982 1842 1985 1868
rect 1990 1822 1993 1848
rect 2006 1802 2009 1858
rect 2014 1852 2017 1868
rect 2022 1862 2025 1868
rect 2078 1862 2081 1868
rect 2102 1862 2105 1908
rect 2174 1872 2177 1878
rect 2070 1852 2073 1858
rect 2054 1842 2057 1848
rect 1998 1762 2001 1788
rect 2002 1748 2006 1751
rect 1966 1732 1969 1738
rect 1974 1712 1977 1748
rect 2030 1742 2033 1768
rect 2066 1758 2070 1761
rect 2086 1752 2089 1798
rect 2102 1792 2105 1848
rect 2142 1831 2145 1850
rect 2122 1788 2126 1791
rect 2110 1742 2113 1778
rect 2118 1752 2121 1758
rect 2134 1752 2137 1828
rect 2018 1738 2022 1741
rect 2066 1738 2070 1741
rect 2098 1738 2102 1741
rect 1982 1732 1985 1738
rect 1982 1672 1985 1688
rect 2006 1672 2009 1738
rect 2026 1728 2030 1731
rect 2054 1722 2057 1728
rect 2026 1688 2030 1691
rect 2026 1678 2030 1681
rect 1994 1668 1998 1671
rect 2042 1668 2046 1671
rect 2006 1662 2009 1668
rect 2054 1662 2057 1698
rect 2062 1682 2065 1728
rect 2094 1712 2097 1738
rect 2134 1722 2137 1738
rect 2150 1732 2153 1808
rect 2190 1762 2193 1878
rect 2230 1852 2233 1858
rect 2222 1752 2225 1808
rect 2158 1742 2161 1748
rect 2102 1712 2105 1718
rect 2134 1692 2137 1718
rect 2142 1702 2145 1728
rect 2150 1692 2153 1728
rect 2106 1688 2110 1691
rect 2062 1662 2065 1668
rect 2078 1662 2081 1678
rect 2126 1672 2129 1678
rect 1990 1642 1993 1658
rect 1858 1528 1862 1531
rect 1854 1472 1857 1528
rect 1870 1491 1873 1538
rect 1918 1532 1921 1538
rect 1880 1503 1882 1507
rect 1886 1503 1889 1507
rect 1893 1503 1896 1507
rect 1958 1492 1961 1598
rect 1966 1542 1969 1618
rect 2094 1592 2097 1668
rect 2110 1642 2113 1668
rect 2118 1652 2121 1658
rect 2126 1591 2129 1668
rect 2190 1602 2193 1718
rect 2198 1702 2201 1738
rect 2210 1728 2214 1731
rect 2230 1692 2233 1758
rect 2246 1742 2249 1758
rect 2254 1752 2257 1918
rect 2294 1902 2297 1948
rect 2262 1772 2265 1888
rect 2294 1882 2297 1888
rect 2274 1878 2278 1881
rect 2302 1872 2305 1948
rect 2326 1942 2329 1948
rect 2314 1938 2318 1941
rect 2314 1928 2318 1931
rect 2314 1898 2321 1901
rect 2318 1872 2321 1898
rect 2350 1892 2353 1938
rect 2366 1892 2369 1908
rect 2298 1868 2302 1871
rect 2286 1732 2289 1868
rect 2306 1858 2310 1861
rect 2310 1752 2313 1848
rect 2326 1842 2329 1848
rect 2334 1802 2337 1868
rect 2358 1862 2361 1878
rect 2366 1862 2369 1868
rect 2350 1842 2353 1848
rect 2374 1822 2377 2008
rect 2384 2003 2386 2007
rect 2390 2003 2393 2007
rect 2397 2003 2400 2007
rect 2398 1952 2401 1988
rect 2382 1932 2385 1948
rect 2406 1942 2409 1958
rect 2414 1952 2417 2068
rect 2450 2058 2454 2061
rect 2422 1952 2425 2058
rect 2430 2032 2433 2038
rect 2446 2002 2449 2048
rect 2470 1992 2473 2038
rect 2430 1962 2433 1968
rect 2478 1962 2481 2088
rect 2530 2078 2534 2081
rect 2570 2078 2577 2081
rect 2550 2072 2553 2078
rect 2574 2072 2577 2078
rect 2586 2068 2590 2071
rect 2602 2068 2606 2071
rect 2542 2062 2545 2068
rect 2566 2062 2569 2068
rect 2614 2062 2617 2208
rect 2622 2192 2625 2218
rect 2638 2162 2641 2178
rect 2586 2058 2590 2061
rect 2486 2052 2489 2058
rect 2506 2048 2510 2051
rect 2510 1962 2513 1978
rect 2438 1952 2441 1958
rect 2446 1952 2449 1958
rect 2450 1938 2454 1941
rect 2466 1938 2470 1941
rect 2422 1932 2425 1938
rect 2418 1918 2422 1921
rect 2470 1892 2473 1918
rect 2478 1892 2481 1938
rect 2446 1882 2449 1888
rect 2426 1878 2430 1881
rect 2430 1872 2433 1878
rect 2466 1868 2470 1871
rect 2390 1852 2393 1858
rect 2384 1803 2386 1807
rect 2390 1803 2393 1807
rect 2397 1803 2400 1807
rect 2366 1732 2369 1738
rect 2238 1701 2241 1718
rect 2238 1698 2249 1701
rect 2230 1682 2233 1688
rect 2246 1672 2249 1698
rect 2314 1678 2318 1681
rect 2330 1668 2334 1671
rect 2298 1658 2302 1661
rect 2122 1588 2129 1591
rect 2070 1560 2073 1579
rect 2090 1548 2094 1551
rect 1982 1542 1985 1548
rect 2038 1542 2041 1548
rect 2022 1522 2025 1528
rect 1870 1488 1878 1491
rect 1942 1482 1945 1488
rect 1870 1462 1873 1468
rect 1906 1458 1910 1461
rect 1838 1422 1841 1428
rect 1814 1408 1825 1411
rect 1822 1392 1825 1408
rect 1838 1362 1841 1418
rect 1810 1358 1814 1361
rect 1846 1352 1849 1448
rect 1830 1342 1833 1348
rect 1846 1342 1849 1348
rect 1746 1338 1753 1341
rect 1738 1328 1742 1331
rect 1750 1312 1753 1338
rect 1790 1338 1798 1341
rect 1718 1292 1721 1298
rect 1758 1292 1761 1338
rect 1790 1292 1793 1338
rect 1738 1288 1742 1291
rect 1706 1268 1710 1271
rect 1726 1261 1729 1278
rect 1778 1268 1782 1271
rect 1726 1258 1734 1261
rect 1638 1232 1641 1258
rect 1734 1252 1737 1258
rect 1750 1252 1753 1268
rect 1806 1262 1809 1288
rect 1758 1242 1761 1248
rect 1718 1222 1721 1228
rect 1614 1168 1625 1171
rect 1622 1162 1625 1168
rect 1618 1148 1622 1151
rect 1606 1142 1609 1148
rect 1638 1142 1641 1168
rect 1646 1152 1649 1218
rect 1654 1202 1657 1218
rect 1590 1138 1601 1141
rect 1590 1122 1593 1128
rect 1582 1118 1590 1121
rect 1574 1092 1577 1118
rect 1598 1092 1601 1138
rect 1606 1122 1609 1138
rect 1618 1128 1622 1131
rect 1634 1128 1638 1131
rect 1630 1092 1633 1118
rect 1474 1078 1481 1081
rect 1462 1072 1465 1078
rect 1442 1068 1446 1071
rect 1470 1062 1473 1068
rect 1478 1062 1481 1078
rect 1494 1062 1497 1078
rect 1502 1062 1505 1068
rect 1494 1052 1497 1058
rect 1474 1048 1478 1051
rect 1510 1042 1513 1058
rect 1526 1052 1529 1078
rect 1622 1072 1625 1078
rect 1586 1068 1590 1071
rect 1622 1062 1625 1068
rect 1638 1062 1641 1068
rect 1662 1062 1665 1178
rect 1686 1142 1689 1198
rect 1734 1172 1737 1238
rect 1742 1192 1745 1218
rect 1806 1192 1809 1258
rect 1762 1188 1766 1191
rect 1670 1122 1673 1128
rect 1670 1072 1673 1078
rect 1678 1072 1681 1088
rect 1710 1072 1713 1088
rect 1718 1062 1721 1148
rect 1690 1058 1694 1061
rect 1534 1052 1537 1058
rect 1550 1002 1553 1018
rect 1334 942 1337 948
rect 1294 892 1297 908
rect 1310 892 1313 908
rect 1310 882 1313 888
rect 1290 878 1294 881
rect 1274 868 1278 871
rect 1230 862 1233 868
rect 1074 858 1078 861
rect 1098 858 1102 861
rect 1202 858 1206 861
rect 1274 858 1278 861
rect 910 822 913 858
rect 1054 831 1057 850
rect 834 768 838 771
rect 774 742 777 748
rect 782 742 785 748
rect 718 682 721 718
rect 734 682 737 728
rect 790 712 793 748
rect 686 622 689 650
rect 718 622 721 668
rect 774 611 777 658
rect 766 608 777 611
rect 766 552 769 608
rect 738 548 742 551
rect 646 532 649 538
rect 630 522 633 528
rect 630 461 633 518
rect 670 482 673 488
rect 622 458 633 461
rect 686 462 689 468
rect 726 462 729 518
rect 758 482 761 518
rect 766 492 769 548
rect 782 462 785 558
rect 558 442 561 458
rect 558 392 561 418
rect 574 402 577 448
rect 594 438 598 441
rect 590 352 593 358
rect 550 322 553 328
rect 462 282 465 288
rect 478 272 481 278
rect 422 262 425 268
rect 518 262 521 308
rect 550 272 553 278
rect 562 258 566 261
rect 318 222 321 250
rect 266 138 270 141
rect 254 122 257 128
rect 254 82 257 118
rect 278 92 281 118
rect 326 62 329 178
rect 334 142 337 248
rect 510 222 513 250
rect 378 218 382 221
rect 344 203 346 207
rect 350 203 353 207
rect 357 203 360 207
rect 446 162 449 188
rect 338 138 342 141
rect 350 62 353 158
rect 494 142 497 208
rect 518 192 521 258
rect 574 252 577 278
rect 582 272 585 308
rect 598 282 601 438
rect 550 152 553 188
rect 510 132 513 138
rect 414 82 417 118
rect 486 82 489 88
rect 502 72 505 78
rect 550 62 553 148
rect 558 62 561 218
rect 590 192 593 198
rect 598 152 601 258
rect 606 142 609 338
rect 614 162 617 168
rect 598 62 601 98
rect 622 92 625 458
rect 630 322 633 328
rect 638 292 641 408
rect 654 352 657 398
rect 726 392 729 458
rect 734 422 737 448
rect 798 442 801 768
rect 818 758 822 761
rect 862 752 865 778
rect 826 748 830 751
rect 814 602 817 618
rect 822 542 825 738
rect 830 692 833 708
rect 848 703 850 707
rect 854 703 857 707
rect 861 703 864 707
rect 838 682 841 698
rect 838 592 841 678
rect 854 562 857 588
rect 850 548 854 551
rect 822 482 825 538
rect 848 503 850 507
rect 854 503 857 507
rect 861 503 864 507
rect 850 468 854 471
rect 822 462 825 468
rect 810 458 814 461
rect 818 448 822 451
rect 750 352 753 388
rect 798 362 801 388
rect 822 352 825 408
rect 657 348 662 351
rect 734 332 737 338
rect 750 332 753 338
rect 674 268 678 271
rect 658 248 662 251
rect 630 162 633 228
rect 638 162 641 218
rect 662 162 665 198
rect 670 182 673 218
rect 694 152 697 258
rect 710 252 713 308
rect 753 268 758 271
rect 750 232 753 268
rect 790 262 793 348
rect 822 332 825 348
rect 838 342 841 468
rect 862 442 865 478
rect 862 362 865 368
rect 870 352 873 658
rect 878 612 881 718
rect 886 692 889 748
rect 958 742 961 828
rect 998 760 1001 779
rect 1030 742 1033 758
rect 1086 752 1089 858
rect 1118 752 1121 818
rect 1126 792 1129 858
rect 1126 772 1129 788
rect 1142 762 1145 818
rect 1166 802 1169 858
rect 1178 848 1182 851
rect 1158 742 1161 778
rect 1206 762 1209 848
rect 1182 752 1185 758
rect 1166 742 1169 748
rect 1174 742 1177 748
rect 1190 742 1193 748
rect 898 738 902 741
rect 1046 732 1049 738
rect 1146 718 1150 721
rect 958 672 961 698
rect 974 682 977 688
rect 1150 682 1153 688
rect 1134 672 1137 678
rect 1014 662 1017 668
rect 1082 658 1086 661
rect 890 648 894 651
rect 910 622 913 648
rect 958 552 961 658
rect 902 542 905 548
rect 918 522 921 528
rect 958 501 961 548
rect 974 522 977 648
rect 1102 631 1105 650
rect 1058 618 1062 621
rect 1054 562 1057 568
rect 1130 558 1134 561
rect 1003 548 1006 551
rect 1014 512 1017 558
rect 1142 552 1145 578
rect 1150 562 1153 568
rect 1158 552 1161 568
rect 1174 552 1177 608
rect 1206 562 1209 758
rect 1222 752 1225 758
rect 1222 732 1225 738
rect 1230 732 1233 738
rect 1230 661 1233 728
rect 1238 712 1241 818
rect 1254 772 1257 788
rect 1254 752 1257 768
rect 1270 732 1273 738
rect 1286 731 1289 878
rect 1302 852 1305 858
rect 1318 762 1321 928
rect 1374 862 1377 948
rect 1398 942 1401 998
rect 1574 992 1577 1038
rect 1450 978 1454 981
rect 1558 952 1561 978
rect 1442 948 1446 951
rect 1570 948 1574 951
rect 1562 938 1566 941
rect 1422 932 1425 938
rect 1454 922 1457 928
rect 1430 902 1433 918
rect 1414 872 1417 878
rect 1430 832 1433 868
rect 1462 831 1465 850
rect 1470 842 1473 918
rect 1326 802 1329 818
rect 1470 812 1473 838
rect 1360 803 1362 807
rect 1366 803 1369 807
rect 1373 803 1376 807
rect 1326 792 1329 798
rect 1282 728 1289 731
rect 1294 712 1297 748
rect 1422 742 1425 778
rect 1334 678 1342 681
rect 1346 678 1350 681
rect 1262 672 1265 678
rect 1230 658 1238 661
rect 1242 658 1246 661
rect 1234 648 1238 651
rect 1254 612 1257 668
rect 1278 662 1281 678
rect 1286 662 1289 678
rect 1318 672 1321 678
rect 1334 672 1337 678
rect 1306 668 1310 671
rect 1346 668 1350 671
rect 1358 662 1361 708
rect 1398 682 1401 688
rect 1406 682 1409 728
rect 1374 672 1377 678
rect 1414 662 1417 668
rect 1454 662 1457 768
rect 1470 762 1473 788
rect 1478 752 1481 858
rect 1494 802 1497 938
rect 1526 902 1529 938
rect 1538 928 1542 931
rect 1506 868 1510 871
rect 1494 732 1497 798
rect 1502 741 1505 868
rect 1534 862 1537 868
rect 1514 858 1518 861
rect 1510 842 1513 848
rect 1510 752 1513 758
rect 1518 752 1521 858
rect 1542 851 1545 918
rect 1550 862 1553 938
rect 1558 872 1561 878
rect 1574 862 1577 948
rect 1582 872 1585 1058
rect 1590 1002 1593 1058
rect 1598 962 1601 1048
rect 1630 1012 1633 1038
rect 1638 1012 1641 1048
rect 1646 1022 1649 1048
rect 1630 962 1633 1008
rect 1686 1002 1689 1018
rect 1594 958 1598 961
rect 1598 942 1601 948
rect 1610 938 1622 941
rect 1626 928 1630 931
rect 1602 888 1606 891
rect 1594 868 1598 871
rect 1614 862 1617 918
rect 1638 882 1641 968
rect 1646 941 1649 978
rect 1682 958 1686 961
rect 1654 952 1657 958
rect 1694 952 1697 1058
rect 1734 1052 1737 1168
rect 1742 1062 1745 1178
rect 1754 1148 1758 1151
rect 1774 1132 1777 1158
rect 1782 1132 1785 1138
rect 1798 1132 1801 1138
rect 1722 1048 1726 1051
rect 1646 938 1654 941
rect 1662 932 1665 938
rect 1686 932 1689 938
rect 1662 862 1665 868
rect 1670 862 1673 918
rect 1678 862 1681 878
rect 1594 858 1598 861
rect 1622 852 1625 858
rect 1646 852 1649 858
rect 1538 848 1545 851
rect 1570 848 1574 851
rect 1526 842 1529 848
rect 1614 822 1617 838
rect 1546 758 1550 761
rect 1578 758 1582 761
rect 1554 748 1558 751
rect 1570 748 1574 751
rect 1502 738 1510 741
rect 1546 738 1550 741
rect 1598 732 1601 758
rect 1614 752 1617 818
rect 1606 732 1609 738
rect 1442 658 1446 661
rect 1310 652 1313 658
rect 1322 648 1326 651
rect 1202 558 1206 561
rect 1214 552 1217 558
rect 1238 551 1241 598
rect 1238 548 1246 551
rect 1030 532 1033 538
rect 1038 532 1041 538
rect 1070 532 1073 538
rect 1078 532 1081 548
rect 1126 542 1129 548
rect 1114 538 1118 541
rect 1158 532 1161 548
rect 1182 542 1185 548
rect 1218 538 1222 541
rect 1166 532 1169 538
rect 1106 528 1110 531
rect 1226 528 1230 531
rect 950 498 961 501
rect 1022 502 1025 518
rect 858 348 862 351
rect 846 342 849 348
rect 874 338 878 341
rect 838 332 841 338
rect 848 303 850 307
rect 854 303 857 307
rect 861 303 864 307
rect 830 282 833 288
rect 846 272 849 278
rect 718 162 721 168
rect 642 148 646 151
rect 698 148 702 151
rect 722 148 726 151
rect 634 138 638 141
rect 690 138 694 141
rect 722 138 726 141
rect 306 58 310 61
rect 586 58 590 61
rect 626 58 630 61
rect 650 58 653 61
rect 262 52 265 58
rect 234 48 238 51
rect 182 22 185 48
rect 182 -19 186 -18
rect 174 -22 186 -19
rect 206 -19 209 18
rect 238 -18 241 48
rect 254 -18 257 48
rect 270 -18 273 38
rect 534 31 537 50
rect 214 -19 218 -18
rect 206 -22 218 -19
rect 238 -22 242 -18
rect 254 -22 258 -18
rect 270 -22 274 -18
rect 286 -19 289 18
rect 294 -19 298 -18
rect 286 -22 298 -19
rect 310 -19 313 18
rect 318 -19 322 -18
rect 310 -22 322 -19
rect 334 -19 337 18
rect 344 3 346 7
rect 350 3 353 7
rect 357 3 360 7
rect 366 -19 370 -18
rect 334 -22 370 -19
rect 374 -19 377 18
rect 382 -19 386 -18
rect 374 -22 386 -19
rect 574 -19 577 18
rect 582 -19 586 -18
rect 574 -22 586 -19
rect 606 -19 610 -18
rect 614 -19 617 18
rect 606 -22 617 -19
rect 630 -19 634 -18
rect 638 -19 641 18
rect 630 -22 641 -19
rect 678 -19 682 -18
rect 686 -19 689 118
rect 710 102 713 138
rect 734 102 737 218
rect 750 162 753 188
rect 734 82 737 88
rect 750 72 753 78
rect 782 12 785 118
rect 790 62 793 258
rect 806 132 809 168
rect 846 152 849 258
rect 886 132 889 478
rect 902 462 905 468
rect 894 362 897 458
rect 910 452 913 498
rect 950 462 953 498
rect 998 482 1001 488
rect 982 472 985 478
rect 918 392 921 448
rect 934 422 937 448
rect 918 362 921 388
rect 926 372 929 378
rect 938 368 942 371
rect 898 348 902 351
rect 910 351 913 358
rect 950 352 953 448
rect 966 372 969 378
rect 1014 362 1017 388
rect 1026 368 1030 371
rect 910 348 921 351
rect 906 338 910 341
rect 918 292 921 348
rect 994 348 998 351
rect 926 342 929 348
rect 1002 338 1006 341
rect 982 332 985 338
rect 934 272 937 328
rect 966 302 969 318
rect 982 312 985 328
rect 950 272 953 278
rect 974 272 977 278
rect 946 258 950 261
rect 962 258 966 261
rect 894 222 897 248
rect 958 222 961 248
rect 974 232 977 268
rect 982 252 985 278
rect 982 182 985 248
rect 990 242 993 258
rect 998 242 1001 298
rect 1014 282 1017 358
rect 1022 342 1025 348
rect 1038 332 1041 458
rect 1054 361 1057 518
rect 1078 492 1081 528
rect 1078 462 1081 488
rect 1094 482 1097 518
rect 1102 492 1105 518
rect 1094 432 1097 468
rect 1118 462 1121 518
rect 1150 502 1153 518
rect 1126 472 1129 478
rect 1134 472 1137 478
rect 1142 472 1145 478
rect 1158 471 1161 528
rect 1150 468 1161 471
rect 1150 462 1153 468
rect 1166 462 1169 518
rect 1174 472 1177 478
rect 1198 472 1201 528
rect 1238 462 1241 548
rect 1262 542 1265 638
rect 1286 592 1289 608
rect 1310 572 1313 648
rect 1334 592 1337 628
rect 1302 552 1305 568
rect 1350 562 1353 648
rect 1362 638 1366 641
rect 1360 603 1362 607
rect 1366 603 1369 607
rect 1373 603 1376 607
rect 1322 548 1326 551
rect 1262 532 1265 538
rect 1278 512 1281 548
rect 1270 462 1273 498
rect 1170 458 1174 461
rect 1234 458 1238 461
rect 1110 402 1113 438
rect 1054 358 1062 361
rect 1046 352 1049 358
rect 1070 352 1073 388
rect 1086 371 1089 388
rect 1082 368 1089 371
rect 1094 352 1097 368
rect 1110 352 1113 388
rect 1146 368 1150 371
rect 1130 348 1134 351
rect 1146 348 1150 351
rect 1046 332 1049 338
rect 1046 322 1049 328
rect 1014 262 1017 268
rect 1022 262 1025 298
rect 1050 288 1054 291
rect 1070 272 1073 308
rect 1078 282 1081 318
rect 1094 282 1097 348
rect 1122 338 1126 341
rect 1102 332 1105 338
rect 1134 332 1137 338
rect 1038 252 1041 268
rect 1046 252 1049 258
rect 1026 238 1030 241
rect 994 218 998 221
rect 1062 212 1065 268
rect 1070 242 1073 268
rect 1110 262 1113 268
rect 1082 258 1086 261
rect 1098 248 1102 251
rect 1106 248 1113 251
rect 1082 218 1086 221
rect 934 160 937 179
rect 982 162 985 168
rect 998 162 1001 168
rect 1022 162 1025 178
rect 1030 172 1033 178
rect 1042 168 1046 171
rect 902 142 905 158
rect 1058 158 1062 161
rect 1030 152 1033 158
rect 986 148 990 151
rect 1002 148 1006 151
rect 1070 151 1073 178
rect 1098 168 1102 171
rect 1110 162 1113 248
rect 1118 242 1121 278
rect 1118 172 1121 238
rect 1134 202 1137 278
rect 1158 262 1161 458
rect 1190 442 1193 458
rect 1166 372 1169 438
rect 1190 342 1193 378
rect 1198 362 1201 368
rect 1206 351 1209 458
rect 1246 432 1249 458
rect 1278 452 1281 458
rect 1286 452 1289 458
rect 1266 438 1270 441
rect 1198 348 1209 351
rect 1182 272 1185 318
rect 1190 312 1193 338
rect 1170 268 1174 271
rect 1182 262 1185 268
rect 1146 258 1150 261
rect 1162 258 1166 261
rect 1198 252 1201 348
rect 1214 302 1217 428
rect 1254 422 1257 428
rect 1246 352 1249 368
rect 1226 348 1233 351
rect 1230 332 1233 348
rect 1246 342 1249 348
rect 1278 332 1281 348
rect 1214 292 1217 298
rect 1214 262 1217 288
rect 1230 262 1233 328
rect 1238 312 1241 318
rect 1294 312 1297 548
rect 1310 542 1313 548
rect 1366 542 1369 548
rect 1342 472 1345 478
rect 1314 458 1318 461
rect 1326 412 1329 468
rect 1350 462 1353 498
rect 1342 442 1345 448
rect 1358 421 1361 518
rect 1366 482 1369 538
rect 1382 472 1385 588
rect 1390 532 1393 558
rect 1390 492 1393 528
rect 1398 502 1401 518
rect 1386 458 1390 461
rect 1350 418 1361 421
rect 1302 382 1305 388
rect 1350 352 1353 418
rect 1360 403 1362 407
rect 1366 403 1369 407
rect 1373 403 1376 407
rect 1318 332 1321 348
rect 1382 341 1385 438
rect 1406 352 1409 658
rect 1462 631 1465 718
rect 1494 692 1497 728
rect 1502 722 1505 728
rect 1542 712 1545 718
rect 1502 692 1505 698
rect 1478 682 1481 688
rect 1494 662 1497 668
rect 1518 662 1521 668
rect 1534 662 1537 698
rect 1566 682 1569 688
rect 1622 682 1625 848
rect 1630 762 1633 848
rect 1678 832 1681 858
rect 1662 822 1665 828
rect 1686 811 1689 928
rect 1694 862 1697 948
rect 1702 932 1705 1048
rect 1758 1032 1761 1078
rect 1710 1012 1713 1018
rect 1710 962 1713 1008
rect 1758 1002 1761 1028
rect 1766 962 1769 1118
rect 1774 1082 1777 1088
rect 1790 1081 1793 1118
rect 1790 1078 1801 1081
rect 1782 1062 1785 1068
rect 1790 992 1793 1068
rect 1798 1062 1801 1078
rect 1778 978 1782 981
rect 1742 952 1745 958
rect 1722 948 1726 951
rect 1766 942 1769 948
rect 1782 942 1785 968
rect 1806 952 1809 1148
rect 1814 1142 1817 1248
rect 1822 1192 1825 1318
rect 1838 1292 1841 1298
rect 1846 1241 1849 1308
rect 1854 1282 1857 1348
rect 1862 1342 1865 1458
rect 1890 1448 1894 1451
rect 1910 1392 1913 1438
rect 1874 1388 1878 1391
rect 1918 1382 1921 1468
rect 1862 1332 1865 1338
rect 1902 1312 1905 1328
rect 1926 1322 1929 1458
rect 1934 1452 1937 1458
rect 2038 1452 2041 1478
rect 2054 1452 2057 1468
rect 2086 1422 2089 1450
rect 2006 1342 2009 1368
rect 2054 1362 2057 1388
rect 1880 1303 1882 1307
rect 1886 1303 1889 1307
rect 1893 1303 1896 1307
rect 1854 1252 1857 1278
rect 1918 1272 1921 1278
rect 1934 1272 1937 1278
rect 1982 1262 1985 1268
rect 1846 1238 1857 1241
rect 1854 1192 1857 1238
rect 1982 1222 1985 1248
rect 1990 1242 1993 1328
rect 2006 1262 2009 1318
rect 2038 1292 2041 1318
rect 2046 1272 2049 1348
rect 2070 1302 2073 1398
rect 2094 1362 2097 1468
rect 2102 1462 2105 1548
rect 2150 1492 2153 1508
rect 2158 1481 2161 1578
rect 2198 1532 2201 1568
rect 2246 1552 2249 1658
rect 2294 1622 2297 1648
rect 2286 1592 2289 1608
rect 2262 1562 2265 1588
rect 2350 1562 2353 1728
rect 2406 1712 2409 1868
rect 2414 1852 2417 1858
rect 2454 1852 2457 1868
rect 2486 1861 2489 1938
rect 2502 1932 2505 1938
rect 2518 1931 2521 2058
rect 2594 2048 2598 2051
rect 2626 2048 2630 2051
rect 2526 1952 2529 1978
rect 2542 1962 2545 1968
rect 2558 1952 2561 2038
rect 2598 1962 2601 1978
rect 2586 1948 2590 1951
rect 2530 1938 2534 1941
rect 2562 1938 2566 1941
rect 2602 1938 2606 1941
rect 2518 1928 2529 1931
rect 2518 1872 2521 1908
rect 2526 1902 2529 1928
rect 2534 1912 2537 1938
rect 2574 1922 2577 1938
rect 2622 1932 2625 2018
rect 2638 1972 2641 2118
rect 2646 2092 2649 2268
rect 2654 2082 2657 2288
rect 2670 2262 2673 2458
rect 2698 2448 2702 2451
rect 2678 2352 2681 2358
rect 2686 2352 2689 2378
rect 2702 2352 2705 2358
rect 2718 2352 2721 2428
rect 2726 2402 2729 2468
rect 2734 2432 2737 2468
rect 2750 2392 2753 2458
rect 2758 2372 2761 2448
rect 2734 2352 2737 2358
rect 2750 2342 2753 2348
rect 2698 2338 2702 2341
rect 2718 2322 2721 2328
rect 2734 2292 2737 2338
rect 2766 2332 2769 2508
rect 2798 2492 2801 2528
rect 2790 2472 2793 2488
rect 2806 2482 2809 2508
rect 2814 2492 2817 2548
rect 2822 2532 2825 2558
rect 2830 2552 2833 2568
rect 2814 2472 2817 2478
rect 2818 2458 2822 2461
rect 2774 2392 2777 2448
rect 2782 2432 2785 2458
rect 2830 2452 2833 2538
rect 2838 2482 2841 2578
rect 2846 2562 2849 2648
rect 2854 2642 2857 2658
rect 2862 2632 2865 2668
rect 2870 2651 2873 2738
rect 2882 2668 2886 2671
rect 2882 2658 2886 2661
rect 2894 2661 2897 2728
rect 2904 2703 2906 2707
rect 2910 2703 2913 2707
rect 2917 2703 2920 2707
rect 2926 2682 2929 2718
rect 2902 2672 2905 2678
rect 2926 2672 2929 2678
rect 2894 2658 2902 2661
rect 2870 2648 2881 2651
rect 2878 2592 2881 2648
rect 2934 2592 2937 2808
rect 2958 2712 2961 2958
rect 2970 2948 2974 2951
rect 2966 2862 2969 2948
rect 2982 2881 2985 2968
rect 2990 2960 2993 2979
rect 3022 2942 3025 3008
rect 3038 2932 3041 3018
rect 3046 3002 3049 3118
rect 3094 3102 3097 3118
rect 3118 3102 3121 3258
rect 3146 3248 3150 3251
rect 3126 3242 3129 3248
rect 3158 3242 3161 3258
rect 3174 3252 3177 3258
rect 3182 3252 3185 3258
rect 3198 3242 3201 3248
rect 3126 3212 3129 3238
rect 3158 3182 3161 3218
rect 3098 3088 3102 3091
rect 3054 3042 3057 3068
rect 3078 3062 3081 3088
rect 3086 3072 3089 3078
rect 3118 3072 3121 3098
rect 3110 3062 3113 3068
rect 3066 3058 3070 3061
rect 3094 3052 3097 3058
rect 3062 3012 3065 3018
rect 2982 2878 2990 2881
rect 2990 2862 2993 2878
rect 2966 2752 2969 2858
rect 3018 2848 3022 2851
rect 3030 2842 3033 2858
rect 3038 2852 3041 2928
rect 3054 2852 3057 2868
rect 3062 2842 3065 2858
rect 3086 2852 3089 2858
rect 3070 2842 3073 2848
rect 3094 2842 3097 2858
rect 3102 2852 3105 2908
rect 3110 2872 3113 3058
rect 3118 2992 3121 3068
rect 3126 3062 3129 3158
rect 3142 3152 3145 3158
rect 3134 3132 3137 3148
rect 3150 3142 3153 3158
rect 3166 3142 3169 3158
rect 3174 3152 3177 3158
rect 3150 3132 3153 3138
rect 3170 3128 3177 3131
rect 3158 3122 3161 3128
rect 3134 3072 3137 3108
rect 3126 3042 3129 3048
rect 3134 2982 3137 3068
rect 3142 3052 3145 3058
rect 3166 3052 3169 3088
rect 3150 3012 3153 3018
rect 3130 2958 3134 2961
rect 3118 2862 3121 2868
rect 3126 2862 3129 2958
rect 3150 2942 3153 2988
rect 3158 2962 3161 2968
rect 3174 2942 3177 3128
rect 3182 3062 3185 3238
rect 3206 3222 3209 3268
rect 3238 3262 3241 3278
rect 3226 3248 3230 3251
rect 3238 3242 3241 3248
rect 3214 3161 3217 3218
rect 3230 3192 3233 3238
rect 3214 3158 3222 3161
rect 3190 3142 3193 3148
rect 3206 3142 3209 3158
rect 3182 2942 3185 2998
rect 3190 2972 3193 3138
rect 3218 3118 3222 3121
rect 3214 3082 3217 3108
rect 3230 3102 3233 3148
rect 3246 3132 3249 3278
rect 3262 3252 3265 3308
rect 3286 3272 3289 3418
rect 3294 3411 3297 3418
rect 3294 3408 3302 3411
rect 3326 3392 3329 3448
rect 3334 3441 3337 3458
rect 3358 3452 3361 3468
rect 3334 3438 3342 3441
rect 3318 3372 3321 3378
rect 3306 3368 3310 3371
rect 3294 3362 3297 3368
rect 3314 3348 3318 3351
rect 3294 3332 3297 3338
rect 3318 3292 3321 3318
rect 3282 3268 3286 3271
rect 3298 3268 3302 3271
rect 3282 3258 3286 3261
rect 3294 3252 3297 3258
rect 3262 3202 3265 3248
rect 3310 3222 3313 3278
rect 3326 3252 3329 3388
rect 3350 3372 3353 3418
rect 3366 3382 3369 3538
rect 3374 3362 3377 3548
rect 3438 3532 3441 3558
rect 3454 3552 3457 3568
rect 3466 3558 3470 3561
rect 3658 3558 3662 3561
rect 3502 3552 3505 3558
rect 3474 3548 3478 3551
rect 3530 3548 3534 3551
rect 3570 3548 3574 3551
rect 3610 3548 3614 3551
rect 3454 3542 3457 3548
rect 3446 3532 3449 3538
rect 3382 3472 3385 3518
rect 3390 3462 3393 3468
rect 3334 3342 3337 3348
rect 3342 3342 3345 3358
rect 3382 3352 3385 3458
rect 3414 3422 3417 3528
rect 3462 3482 3465 3548
rect 3478 3542 3481 3548
rect 3478 3522 3481 3528
rect 3510 3522 3513 3528
rect 3518 3492 3521 3528
rect 3514 3478 3518 3481
rect 3430 3462 3433 3478
rect 3438 3462 3441 3468
rect 3462 3432 3465 3468
rect 3478 3462 3481 3468
rect 3494 3442 3497 3448
rect 3362 3348 3366 3351
rect 3334 3270 3337 3298
rect 3342 3292 3345 3338
rect 3350 3332 3353 3338
rect 3342 3272 3345 3278
rect 3350 3272 3353 3278
rect 3358 3262 3361 3348
rect 3382 3332 3385 3338
rect 3378 3318 3382 3321
rect 3398 3312 3401 3418
rect 3454 3412 3457 3418
rect 3408 3403 3410 3407
rect 3414 3403 3417 3407
rect 3421 3403 3424 3407
rect 3486 3392 3489 3418
rect 3502 3402 3505 3448
rect 3518 3432 3521 3468
rect 3526 3462 3529 3548
rect 3550 3542 3553 3548
rect 3542 3502 3545 3538
rect 3646 3532 3649 3548
rect 3662 3542 3665 3548
rect 3566 3512 3569 3518
rect 3566 3462 3569 3508
rect 3582 3492 3585 3518
rect 3590 3502 3593 3528
rect 3598 3522 3601 3528
rect 3606 3482 3609 3518
rect 3546 3458 3550 3461
rect 3582 3452 3585 3468
rect 3622 3462 3625 3468
rect 3530 3438 3534 3441
rect 3542 3432 3545 3448
rect 3590 3442 3593 3448
rect 3562 3438 3566 3441
rect 3546 3418 3550 3421
rect 3574 3412 3577 3418
rect 3430 3372 3433 3388
rect 3478 3362 3481 3388
rect 3426 3358 3430 3361
rect 3406 3342 3409 3358
rect 3438 3322 3441 3348
rect 3486 3342 3489 3348
rect 3398 3262 3401 3278
rect 3406 3272 3409 3318
rect 3406 3262 3409 3268
rect 3370 3258 3374 3261
rect 3426 3258 3430 3261
rect 3398 3252 3401 3258
rect 3386 3248 3390 3251
rect 3438 3242 3441 3248
rect 3262 3172 3265 3178
rect 3254 3132 3257 3138
rect 3202 3078 3206 3081
rect 3238 3072 3241 3118
rect 3210 3068 3214 3071
rect 3230 3052 3233 3058
rect 3238 3052 3241 3058
rect 3230 2952 3233 2968
rect 3238 2962 3241 3038
rect 3230 2942 3233 2948
rect 3150 2922 3153 2938
rect 3174 2932 3177 2938
rect 3238 2932 3241 2958
rect 3246 2931 3249 3128
rect 3262 3122 3265 3148
rect 3254 3072 3257 3088
rect 3270 3081 3273 3208
rect 3278 3162 3281 3178
rect 3318 3162 3321 3218
rect 3350 3182 3353 3218
rect 3286 3132 3289 3148
rect 3302 3132 3305 3148
rect 3318 3132 3321 3148
rect 3326 3142 3329 3148
rect 3294 3081 3297 3118
rect 3270 3078 3281 3081
rect 3254 3062 3257 3068
rect 3262 3062 3265 3068
rect 3270 3022 3273 3068
rect 3278 3062 3281 3078
rect 3286 3078 3297 3081
rect 3286 3051 3289 3078
rect 3310 3071 3313 3118
rect 3306 3068 3313 3071
rect 3294 3062 3297 3068
rect 3334 3062 3337 3158
rect 3342 3132 3345 3158
rect 3358 3142 3361 3148
rect 3366 3141 3369 3198
rect 3374 3152 3377 3218
rect 3408 3203 3410 3207
rect 3414 3203 3417 3207
rect 3421 3203 3424 3207
rect 3430 3162 3433 3218
rect 3386 3158 3390 3161
rect 3446 3161 3449 3318
rect 3454 3262 3457 3338
rect 3462 3322 3465 3338
rect 3490 3328 3494 3331
rect 3478 3282 3481 3288
rect 3502 3282 3505 3398
rect 3598 3392 3601 3438
rect 3606 3422 3609 3458
rect 3518 3358 3526 3361
rect 3562 3358 3566 3361
rect 3510 3342 3513 3358
rect 3518 3352 3521 3358
rect 3554 3348 3558 3351
rect 3526 3342 3529 3348
rect 3466 3278 3470 3281
rect 3490 3258 3494 3261
rect 3442 3158 3449 3161
rect 3398 3142 3401 3158
rect 3470 3152 3473 3258
rect 3502 3242 3505 3278
rect 3510 3262 3513 3338
rect 3530 3328 3534 3331
rect 3518 3272 3521 3278
rect 3526 3252 3529 3258
rect 3534 3252 3537 3298
rect 3542 3292 3545 3318
rect 3550 3272 3553 3338
rect 3546 3258 3550 3261
rect 3542 3232 3545 3248
rect 3438 3142 3441 3148
rect 3446 3142 3449 3148
rect 3486 3142 3489 3218
rect 3502 3162 3505 3218
rect 3550 3211 3553 3238
rect 3558 3221 3561 3348
rect 3582 3342 3585 3368
rect 3590 3342 3593 3358
rect 3598 3352 3601 3368
rect 3606 3352 3609 3418
rect 3614 3382 3617 3448
rect 3630 3442 3633 3518
rect 3646 3492 3649 3498
rect 3670 3472 3673 3518
rect 3686 3492 3689 3568
rect 3710 3532 3713 3548
rect 3734 3532 3737 3540
rect 3742 3532 3745 3538
rect 3694 3492 3697 3518
rect 3662 3442 3665 3468
rect 3670 3442 3673 3458
rect 3702 3452 3705 3458
rect 3682 3448 3686 3451
rect 3630 3402 3633 3418
rect 3622 3352 3625 3358
rect 3630 3342 3633 3368
rect 3654 3332 3657 3428
rect 3694 3402 3697 3448
rect 3702 3422 3705 3428
rect 3710 3411 3713 3438
rect 3702 3408 3713 3411
rect 3670 3352 3673 3378
rect 3682 3348 3686 3351
rect 3670 3332 3673 3348
rect 3678 3338 3686 3341
rect 3638 3322 3641 3328
rect 3566 3231 3569 3318
rect 3614 3301 3617 3318
rect 3646 3302 3649 3328
rect 3662 3322 3665 3328
rect 3614 3298 3625 3301
rect 3578 3258 3582 3261
rect 3606 3252 3609 3268
rect 3614 3262 3617 3288
rect 3622 3281 3625 3298
rect 3638 3282 3641 3288
rect 3622 3278 3630 3281
rect 3622 3252 3625 3278
rect 3642 3268 3646 3271
rect 3650 3258 3654 3261
rect 3590 3242 3593 3248
rect 3578 3238 3582 3241
rect 3566 3228 3577 3231
rect 3558 3218 3569 3221
rect 3550 3208 3561 3211
rect 3558 3192 3561 3208
rect 3550 3172 3553 3178
rect 3566 3172 3569 3218
rect 3546 3168 3550 3171
rect 3566 3162 3569 3168
rect 3366 3138 3374 3141
rect 3410 3138 3414 3141
rect 3390 3132 3393 3138
rect 3350 3082 3353 3088
rect 3374 3072 3377 3098
rect 3398 3092 3401 3128
rect 3302 3051 3305 3058
rect 3366 3052 3369 3058
rect 3286 3048 3305 3051
rect 3254 2972 3257 3018
rect 3294 3012 3297 3038
rect 3326 3022 3329 3048
rect 3382 3042 3385 3058
rect 3398 3042 3401 3048
rect 3406 3022 3409 3068
rect 3414 3022 3417 3138
rect 3438 3132 3441 3138
rect 3478 3122 3481 3138
rect 3486 3132 3489 3138
rect 3502 3132 3505 3148
rect 3518 3132 3521 3138
rect 3534 3132 3537 3138
rect 3430 3062 3433 3078
rect 3462 3071 3465 3118
rect 3478 3081 3481 3118
rect 3478 3078 3486 3081
rect 3458 3068 3465 3071
rect 3510 3072 3513 3078
rect 3518 3062 3521 3128
rect 3526 3092 3529 3118
rect 3466 3058 3470 3061
rect 3482 3058 3486 3061
rect 3498 3058 3502 3061
rect 3310 3012 3313 3018
rect 3408 3003 3410 3007
rect 3414 3003 3417 3007
rect 3421 3003 3424 3007
rect 3334 2972 3337 2988
rect 3342 2972 3345 2978
rect 3274 2968 3278 2971
rect 3354 2968 3361 2971
rect 3254 2942 3257 2968
rect 3318 2962 3321 2968
rect 3350 2962 3353 2968
rect 3290 2958 3294 2961
rect 3342 2952 3345 2958
rect 3330 2948 3334 2951
rect 3262 2932 3265 2948
rect 3246 2928 3257 2931
rect 3142 2852 3145 2918
rect 3166 2892 3169 2918
rect 3214 2902 3217 2918
rect 3246 2892 3249 2918
rect 3150 2872 3153 2878
rect 3206 2872 3209 2878
rect 3254 2872 3257 2928
rect 3270 2892 3273 2938
rect 3286 2932 3289 2948
rect 3302 2942 3305 2948
rect 3318 2942 3321 2948
rect 3358 2932 3361 2968
rect 3414 2962 3417 2978
rect 3386 2948 3390 2951
rect 3374 2942 3377 2948
rect 3262 2882 3265 2888
rect 3198 2862 3201 2868
rect 3150 2852 3153 2858
rect 3102 2842 3105 2848
rect 2994 2838 2998 2841
rect 2998 2792 3001 2838
rect 3038 2832 3041 2838
rect 3070 2832 3073 2838
rect 3234 2828 3238 2831
rect 3046 2801 3049 2818
rect 3046 2798 3057 2801
rect 3022 2742 3025 2748
rect 3006 2732 3009 2738
rect 3054 2702 3057 2798
rect 3070 2762 3073 2788
rect 3078 2772 3081 2818
rect 3078 2752 3081 2758
rect 3046 2682 3049 2688
rect 2946 2668 2950 2671
rect 3030 2662 3033 2668
rect 3086 2662 3089 2748
rect 2942 2592 2945 2658
rect 2962 2648 2966 2651
rect 3094 2652 3097 2818
rect 3126 2802 3129 2818
rect 3126 2760 3129 2779
rect 3106 2748 3110 2751
rect 3158 2742 3161 2798
rect 3254 2792 3257 2868
rect 3262 2862 3265 2878
rect 3278 2872 3281 2918
rect 3310 2882 3313 2918
rect 3358 2892 3361 2928
rect 3390 2922 3393 2938
rect 3370 2918 3374 2921
rect 3370 2878 3374 2881
rect 3310 2872 3313 2878
rect 3298 2848 3302 2851
rect 3318 2832 3321 2878
rect 3334 2862 3337 2868
rect 3330 2848 3334 2851
rect 3342 2842 3345 2848
rect 3358 2832 3361 2858
rect 3174 2722 3177 2728
rect 3142 2652 3145 2698
rect 3166 2682 3169 2698
rect 3238 2682 3241 2788
rect 3294 2762 3297 2768
rect 3270 2752 3273 2758
rect 3262 2742 3265 2748
rect 3278 2741 3281 2748
rect 3274 2738 3281 2741
rect 3302 2742 3305 2828
rect 3366 2822 3369 2828
rect 3350 2772 3353 2818
rect 3358 2752 3361 2758
rect 3374 2752 3377 2878
rect 3382 2872 3385 2918
rect 3386 2858 3390 2861
rect 3398 2832 3401 2948
rect 3422 2882 3425 2938
rect 3422 2872 3425 2878
rect 3406 2832 3409 2848
rect 3382 2752 3385 2768
rect 3358 2732 3361 2748
rect 3374 2732 3377 2748
rect 3390 2742 3393 2818
rect 3408 2803 3410 2807
rect 3414 2803 3417 2807
rect 3421 2803 3424 2807
rect 3430 2802 3433 3048
rect 3438 2792 3441 3058
rect 3450 3048 3454 3051
rect 3462 3042 3465 3048
rect 3446 2952 3449 2988
rect 3454 2972 3457 3018
rect 3478 3002 3481 3048
rect 3510 3022 3513 3058
rect 3530 3048 3534 3051
rect 3518 3042 3521 3048
rect 3550 3042 3553 3158
rect 3574 3152 3577 3228
rect 3562 3148 3566 3151
rect 3574 3142 3577 3148
rect 3558 3062 3561 3118
rect 3582 3062 3585 3218
rect 3590 3162 3593 3238
rect 3598 3162 3601 3218
rect 3614 3162 3617 3238
rect 3622 3158 3630 3161
rect 3614 3152 3617 3158
rect 3622 3152 3625 3158
rect 3654 3152 3657 3258
rect 3662 3252 3665 3298
rect 3678 3262 3681 3308
rect 3694 3282 3697 3318
rect 3686 3272 3689 3278
rect 3702 3222 3705 3408
rect 3718 3382 3721 3518
rect 3726 3472 3729 3478
rect 3742 3472 3745 3478
rect 3758 3472 3761 3498
rect 3726 3372 3729 3418
rect 3722 3358 3726 3361
rect 3714 3338 3718 3341
rect 3714 3328 3718 3331
rect 3734 3321 3737 3398
rect 3742 3372 3745 3468
rect 3750 3412 3753 3458
rect 3774 3442 3777 3448
rect 3754 3408 3761 3411
rect 3750 3342 3753 3358
rect 3758 3352 3761 3408
rect 3742 3332 3745 3338
rect 3758 3332 3761 3338
rect 3734 3318 3745 3321
rect 3726 3302 3729 3318
rect 3734 3272 3737 3308
rect 3742 3292 3745 3318
rect 3766 3282 3769 3418
rect 3746 3278 3750 3281
rect 3774 3262 3777 3368
rect 3722 3258 3726 3261
rect 3710 3252 3713 3258
rect 3766 3252 3769 3258
rect 3722 3248 3726 3251
rect 3718 3242 3721 3248
rect 3678 3192 3681 3218
rect 3718 3192 3721 3218
rect 3602 3138 3606 3141
rect 3590 3122 3593 3128
rect 3586 3048 3590 3051
rect 3462 2982 3465 2988
rect 3518 2982 3521 3028
rect 3502 2962 3505 2968
rect 3470 2942 3473 2948
rect 3518 2942 3521 2978
rect 3526 2942 3529 3018
rect 3538 2958 3542 2961
rect 3558 2961 3561 3018
rect 3550 2958 3561 2961
rect 3566 3002 3569 3048
rect 3586 3038 3590 3041
rect 3542 2942 3545 2948
rect 3550 2942 3553 2958
rect 3526 2932 3529 2938
rect 3454 2892 3457 2928
rect 3462 2852 3465 2928
rect 3470 2872 3473 2888
rect 3518 2872 3521 2878
rect 3526 2872 3529 2898
rect 3550 2871 3553 2938
rect 3558 2902 3561 2940
rect 3566 2922 3569 2998
rect 3574 2932 3577 3018
rect 3614 2992 3617 3148
rect 3654 3142 3657 3148
rect 3662 3142 3665 3148
rect 3686 3142 3689 3168
rect 3702 3162 3705 3178
rect 3710 3162 3713 3168
rect 3718 3152 3721 3168
rect 3726 3162 3729 3168
rect 3742 3132 3745 3138
rect 3750 3132 3753 3218
rect 3650 3128 3654 3131
rect 3638 3091 3641 3118
rect 3638 3088 3649 3091
rect 3634 3078 3638 3081
rect 3646 3071 3649 3088
rect 3654 3082 3657 3128
rect 3678 3122 3681 3128
rect 3670 3072 3673 3118
rect 3702 3092 3705 3118
rect 3706 3078 3710 3081
rect 3642 3068 3649 3071
rect 3658 3068 3662 3071
rect 3678 3062 3681 3078
rect 3718 3072 3721 3088
rect 3726 3062 3729 3118
rect 3750 3102 3753 3128
rect 3766 3082 3769 3228
rect 3738 3068 3742 3071
rect 3626 3058 3630 3061
rect 3746 3058 3750 3061
rect 3582 2952 3585 2968
rect 3566 2892 3569 2918
rect 3574 2882 3577 2918
rect 3582 2881 3585 2948
rect 3590 2942 3593 2978
rect 3622 2962 3625 3018
rect 3646 2952 3649 3058
rect 3662 3052 3665 3058
rect 3694 3052 3697 3058
rect 3738 3048 3742 3051
rect 3678 2971 3681 3018
rect 3674 2968 3681 2971
rect 3654 2952 3657 2958
rect 3686 2952 3689 3008
rect 3610 2948 3614 2951
rect 3666 2948 3670 2951
rect 3662 2942 3665 2948
rect 3626 2938 3630 2941
rect 3642 2938 3646 2941
rect 3582 2878 3593 2881
rect 3542 2868 3553 2871
rect 3578 2868 3582 2871
rect 3542 2852 3545 2868
rect 3590 2862 3593 2878
rect 3458 2848 3462 2851
rect 3438 2772 3441 2778
rect 3446 2742 3449 2838
rect 3454 2762 3457 2848
rect 3550 2832 3553 2858
rect 3598 2851 3601 2918
rect 3606 2882 3609 2928
rect 3634 2868 3638 2871
rect 3646 2871 3649 2918
rect 3654 2882 3657 2938
rect 3702 2932 3705 3038
rect 3734 2951 3737 2958
rect 3730 2948 3737 2951
rect 3758 2952 3761 3018
rect 3770 2948 3774 2951
rect 3694 2922 3697 2928
rect 3662 2912 3665 2918
rect 3646 2868 3654 2871
rect 3614 2862 3617 2868
rect 3598 2848 3606 2851
rect 3590 2842 3593 2848
rect 3498 2818 3502 2821
rect 3454 2752 3457 2758
rect 3470 2742 3473 2758
rect 3494 2742 3497 2798
rect 3534 2772 3537 2818
rect 3542 2762 3545 2818
rect 3502 2752 3505 2758
rect 3518 2742 3521 2758
rect 3566 2752 3569 2778
rect 3598 2762 3601 2778
rect 3630 2752 3633 2828
rect 3662 2762 3665 2878
rect 3670 2862 3673 2888
rect 3710 2871 3713 2918
rect 3726 2882 3729 2948
rect 3738 2938 3742 2941
rect 3734 2882 3737 2928
rect 3710 2868 3718 2871
rect 3686 2862 3689 2868
rect 3742 2862 3745 2938
rect 3758 2932 3761 2938
rect 3750 2922 3753 2928
rect 3766 2892 3769 2918
rect 3762 2878 3766 2881
rect 3694 2762 3697 2848
rect 3726 2772 3729 2778
rect 3750 2772 3753 2818
rect 3714 2768 3718 2771
rect 3690 2758 3694 2761
rect 3750 2758 3758 2761
rect 3554 2748 3558 2751
rect 3618 2748 3622 2751
rect 3566 2742 3569 2748
rect 3426 2738 3430 2741
rect 3498 2738 3505 2741
rect 3410 2728 3414 2731
rect 3402 2718 3406 2721
rect 3294 2712 3297 2718
rect 3262 2692 3265 2708
rect 3178 2678 3182 2681
rect 3166 2672 3169 2678
rect 3262 2672 3265 2688
rect 3326 2682 3329 2718
rect 3334 2712 3337 2718
rect 3486 2702 3489 2718
rect 3350 2682 3353 2698
rect 3486 2682 3489 2688
rect 3290 2678 3294 2681
rect 3454 2678 3462 2681
rect 3194 2668 3198 2671
rect 3274 2668 3278 2671
rect 3290 2668 3294 2671
rect 3158 2662 3161 2668
rect 3194 2658 3198 2661
rect 2998 2622 3001 2650
rect 3122 2638 3126 2641
rect 3190 2632 3193 2658
rect 3202 2648 3206 2651
rect 2990 2592 2993 2598
rect 2854 2562 2857 2588
rect 2862 2562 2865 2568
rect 2958 2562 2961 2578
rect 2850 2558 2854 2561
rect 2870 2558 2889 2561
rect 2870 2551 2873 2558
rect 2866 2548 2873 2551
rect 2886 2551 2889 2558
rect 2974 2552 2977 2558
rect 2886 2548 2910 2551
rect 2854 2492 2857 2528
rect 2878 2511 2881 2548
rect 2982 2542 2985 2548
rect 2998 2542 3001 2608
rect 3034 2558 3038 2561
rect 3034 2548 3038 2551
rect 2898 2538 2902 2541
rect 2930 2538 2937 2541
rect 2886 2532 2889 2538
rect 2894 2518 2902 2521
rect 2878 2508 2886 2511
rect 2894 2502 2897 2518
rect 2904 2503 2906 2507
rect 2910 2503 2913 2507
rect 2917 2503 2920 2507
rect 2894 2492 2897 2498
rect 2934 2492 2937 2538
rect 3006 2531 3009 2548
rect 3046 2542 3049 2578
rect 3062 2542 3065 2548
rect 3070 2542 3073 2568
rect 3086 2562 3089 2578
rect 3094 2542 3097 2618
rect 3110 2562 3113 2578
rect 3158 2552 3161 2618
rect 3174 2562 3177 2618
rect 3182 2562 3185 2568
rect 3170 2548 3174 2551
rect 2998 2528 3009 2531
rect 3066 2528 3070 2531
rect 2838 2472 2841 2478
rect 2846 2462 2849 2478
rect 2862 2462 2865 2468
rect 2870 2462 2873 2488
rect 2882 2468 2886 2471
rect 2894 2462 2897 2488
rect 2926 2472 2929 2478
rect 2942 2472 2945 2528
rect 2986 2478 2990 2481
rect 2958 2472 2961 2478
rect 2998 2472 3001 2528
rect 3014 2482 3017 2528
rect 3010 2468 3014 2471
rect 2902 2462 2905 2468
rect 2798 2352 2801 2438
rect 2814 2392 2817 2398
rect 2838 2392 2841 2418
rect 2794 2338 2798 2341
rect 2806 2332 2809 2338
rect 2810 2328 2822 2331
rect 2774 2322 2777 2328
rect 2734 2272 2737 2278
rect 2774 2272 2777 2318
rect 2830 2302 2833 2388
rect 2846 2352 2849 2458
rect 2870 2352 2873 2388
rect 2878 2352 2881 2448
rect 2822 2272 2825 2278
rect 2830 2272 2833 2298
rect 2718 2262 2721 2268
rect 2778 2258 2782 2261
rect 2686 2231 2689 2250
rect 2814 2222 2817 2248
rect 2758 2162 2761 2178
rect 2674 2158 2678 2161
rect 2698 2158 2702 2161
rect 2722 2158 2729 2161
rect 2662 2152 2665 2158
rect 2726 2152 2729 2158
rect 2682 2148 2686 2151
rect 2746 2148 2750 2151
rect 2718 2142 2721 2148
rect 2662 2092 2665 2138
rect 2670 2112 2673 2118
rect 2654 2072 2657 2078
rect 2662 2062 2665 2068
rect 2670 2062 2673 2098
rect 2686 2082 2689 2118
rect 2694 2102 2697 2138
rect 2726 2132 2729 2138
rect 2734 2112 2737 2138
rect 2734 2092 2737 2098
rect 2726 2072 2729 2078
rect 2758 2072 2761 2158
rect 2774 2142 2777 2188
rect 2806 2162 2809 2188
rect 2814 2172 2817 2218
rect 2838 2182 2841 2348
rect 2862 2342 2865 2348
rect 2850 2338 2854 2341
rect 2874 2338 2878 2341
rect 2862 2292 2865 2298
rect 2894 2292 2897 2368
rect 2904 2303 2906 2307
rect 2910 2303 2913 2307
rect 2917 2303 2920 2307
rect 2942 2292 2945 2468
rect 2954 2458 2958 2461
rect 2970 2458 2974 2461
rect 2982 2452 2985 2468
rect 2998 2462 3001 2468
rect 2990 2452 2993 2458
rect 2998 2362 3001 2458
rect 3022 2452 3025 2478
rect 3030 2462 3033 2518
rect 3086 2482 3089 2518
rect 3094 2482 3097 2518
rect 3062 2472 3065 2478
rect 3070 2472 3073 2478
rect 3030 2372 3033 2418
rect 3038 2351 3041 2438
rect 3058 2428 3062 2431
rect 3046 2362 3049 2388
rect 3038 2348 3049 2351
rect 2998 2342 3001 2348
rect 3030 2342 3033 2348
rect 2982 2332 2985 2338
rect 3006 2292 3009 2308
rect 2954 2288 2958 2291
rect 2942 2282 2945 2288
rect 2886 2272 2889 2278
rect 2950 2272 2953 2288
rect 2974 2282 2977 2288
rect 3038 2282 3041 2318
rect 3046 2292 3049 2348
rect 3030 2272 3033 2278
rect 3038 2272 3041 2278
rect 3062 2272 3065 2358
rect 3070 2352 3073 2418
rect 3078 2372 3081 2418
rect 3086 2362 3089 2448
rect 3102 2431 3105 2528
rect 3118 2522 3121 2548
rect 3166 2538 3174 2541
rect 3190 2538 3198 2541
rect 3154 2528 3158 2531
rect 3134 2492 3137 2518
rect 3142 2512 3145 2518
rect 3166 2492 3169 2538
rect 3110 2462 3113 2468
rect 3118 2462 3121 2488
rect 3146 2478 3150 2481
rect 3146 2468 3150 2471
rect 3094 2428 3105 2431
rect 3070 2302 3073 2348
rect 3078 2342 3081 2358
rect 3094 2332 3097 2428
rect 3126 2422 3129 2468
rect 3174 2462 3177 2498
rect 3190 2492 3193 2538
rect 3206 2481 3209 2588
rect 3214 2582 3217 2668
rect 3222 2662 3225 2668
rect 3230 2652 3233 2668
rect 3326 2662 3329 2668
rect 3258 2658 3265 2661
rect 3230 2622 3233 2648
rect 3214 2562 3217 2578
rect 3222 2562 3225 2618
rect 3254 2612 3257 2618
rect 3254 2562 3257 2578
rect 3262 2562 3265 2658
rect 3238 2542 3241 2558
rect 3262 2551 3265 2558
rect 3254 2548 3265 2551
rect 3286 2551 3289 2618
rect 3326 2572 3329 2658
rect 3318 2562 3321 2568
rect 3286 2548 3294 2551
rect 3226 2538 3230 2541
rect 3222 2492 3225 2518
rect 3238 2488 3246 2491
rect 3202 2478 3209 2481
rect 3230 2482 3233 2488
rect 3238 2482 3241 2488
rect 3242 2468 3246 2471
rect 3166 2442 3169 2448
rect 3182 2442 3185 2468
rect 3106 2418 3110 2421
rect 3118 2352 3121 2358
rect 3134 2342 3137 2438
rect 3166 2422 3169 2438
rect 3206 2382 3209 2458
rect 3214 2442 3217 2468
rect 3254 2462 3257 2548
rect 3278 2538 3286 2541
rect 3262 2522 3265 2538
rect 3278 2492 3281 2538
rect 3294 2531 3297 2538
rect 3290 2528 3297 2531
rect 3326 2532 3329 2548
rect 3334 2531 3337 2648
rect 3342 2642 3345 2648
rect 3350 2562 3353 2658
rect 3342 2552 3345 2558
rect 3366 2552 3369 2658
rect 3382 2652 3385 2658
rect 3374 2552 3377 2608
rect 3366 2542 3369 2548
rect 3334 2528 3342 2531
rect 3262 2472 3265 2488
rect 3230 2362 3233 2368
rect 3154 2358 3158 2361
rect 3262 2352 3265 2388
rect 3170 2348 3174 2351
rect 3210 2348 3214 2351
rect 3122 2338 3126 2341
rect 3170 2338 3174 2341
rect 3194 2338 3198 2341
rect 3250 2338 3254 2341
rect 3078 2282 3081 2318
rect 2994 2268 2998 2271
rect 3050 2268 3054 2271
rect 2826 2148 2830 2151
rect 2790 2142 2793 2148
rect 2842 2138 2846 2141
rect 2782 2132 2785 2138
rect 2822 2132 2825 2138
rect 2766 2122 2769 2128
rect 2854 2102 2857 2258
rect 2866 2188 2870 2191
rect 2822 2082 2825 2088
rect 2806 2072 2809 2078
rect 2706 2058 2710 2061
rect 2662 2052 2665 2058
rect 2694 2042 2697 2048
rect 2674 2038 2678 2041
rect 2662 1962 2665 2038
rect 2718 2002 2721 2068
rect 2862 2062 2865 2148
rect 2878 2131 2881 2258
rect 2902 2192 2905 2258
rect 2934 2252 2937 2268
rect 3022 2262 3025 2268
rect 2962 2258 2966 2261
rect 2994 2258 2998 2261
rect 2982 2252 2985 2258
rect 3002 2248 3006 2251
rect 2910 2212 2913 2218
rect 3014 2162 3017 2188
rect 3022 2152 3025 2188
rect 2906 2148 2910 2151
rect 2950 2132 2953 2138
rect 2966 2132 2969 2138
rect 3030 2132 3033 2268
rect 3102 2262 3105 2318
rect 3134 2312 3137 2338
rect 3182 2332 3185 2338
rect 3158 2322 3161 2328
rect 3110 2272 3113 2278
rect 3150 2272 3153 2318
rect 3050 2258 3054 2261
rect 3038 2192 3041 2258
rect 3102 2242 3105 2248
rect 3070 2192 3073 2218
rect 3102 2142 3105 2198
rect 3110 2162 3113 2258
rect 3118 2252 3121 2258
rect 3126 2252 3129 2258
rect 3134 2242 3137 2248
rect 3126 2172 3129 2218
rect 3150 2192 3153 2258
rect 3166 2252 3169 2258
rect 3122 2158 3126 2161
rect 3110 2142 3113 2148
rect 3050 2138 3054 2141
rect 3082 2138 3086 2141
rect 2878 2128 2886 2131
rect 2904 2103 2906 2107
rect 2910 2103 2913 2107
rect 2917 2103 2920 2107
rect 2990 2092 2993 2098
rect 2966 2082 2969 2088
rect 2950 2072 2953 2078
rect 2954 2058 2958 2061
rect 2758 2022 2761 2048
rect 2806 2022 2809 2058
rect 2898 2028 2902 2031
rect 2742 2002 2745 2018
rect 2718 1972 2721 1998
rect 2702 1958 2734 1961
rect 2650 1938 2654 1941
rect 2686 1932 2689 1938
rect 2694 1922 2697 1958
rect 2702 1942 2705 1958
rect 2710 1942 2713 1948
rect 2718 1942 2721 1948
rect 2530 1898 2537 1901
rect 2534 1872 2537 1898
rect 2506 1868 2510 1871
rect 2542 1862 2545 1918
rect 2638 1901 2641 1918
rect 2726 1902 2729 1938
rect 2734 1922 2737 1948
rect 2638 1898 2649 1901
rect 2646 1872 2649 1898
rect 2662 1872 2665 1878
rect 2474 1858 2489 1861
rect 2498 1858 2502 1861
rect 2522 1858 2526 1861
rect 2486 1822 2489 1848
rect 2414 1762 2417 1788
rect 2458 1758 2462 1761
rect 2474 1758 2486 1761
rect 2502 1752 2505 1818
rect 2514 1758 2518 1761
rect 2370 1688 2374 1691
rect 2362 1678 2366 1681
rect 2414 1662 2417 1748
rect 2470 1702 2473 1748
rect 2486 1742 2489 1748
rect 2514 1738 2518 1741
rect 2478 1732 2481 1738
rect 2358 1592 2361 1618
rect 2384 1603 2386 1607
rect 2390 1603 2393 1607
rect 2397 1603 2400 1607
rect 2454 1562 2457 1678
rect 2470 1672 2473 1688
rect 2502 1631 2505 1650
rect 2502 1562 2505 1588
rect 2214 1542 2217 1548
rect 2246 1532 2249 1548
rect 2294 1532 2297 1538
rect 2150 1478 2161 1481
rect 2078 1342 2081 1348
rect 2070 1292 2073 1298
rect 2046 1262 2049 1268
rect 2102 1262 2105 1458
rect 2126 1442 2129 1468
rect 2134 1372 2137 1418
rect 2118 1362 2121 1368
rect 2134 1352 2137 1358
rect 2126 1332 2129 1338
rect 2150 1282 2153 1478
rect 2230 1462 2233 1478
rect 2246 1472 2249 1498
rect 2278 1462 2281 1528
rect 2190 1402 2193 1458
rect 2222 1398 2230 1401
rect 2162 1358 2166 1361
rect 2162 1338 2166 1341
rect 2182 1332 2185 1348
rect 2190 1342 2193 1368
rect 2198 1342 2201 1348
rect 2182 1312 2185 1328
rect 2018 1258 2022 1261
rect 2106 1258 2110 1261
rect 2006 1232 2009 1258
rect 1902 1162 1905 1208
rect 1938 1188 1942 1191
rect 1922 1178 1926 1181
rect 1862 1152 1865 1158
rect 1818 1138 1822 1141
rect 1862 1132 1865 1138
rect 1878 1121 1881 1138
rect 1870 1118 1881 1121
rect 1902 1122 1905 1158
rect 1918 1152 1921 1158
rect 1822 1032 1825 1118
rect 1870 1112 1873 1118
rect 1926 1112 1929 1138
rect 2022 1132 2025 1218
rect 2038 1152 2041 1218
rect 2054 1202 2057 1258
rect 2070 1160 2073 1179
rect 2086 1152 2089 1258
rect 2038 1122 2041 1138
rect 1880 1103 1882 1107
rect 1886 1103 1889 1107
rect 1893 1103 1896 1107
rect 1942 1102 1945 1118
rect 1830 1062 1833 1098
rect 1998 1092 2001 1108
rect 1894 1082 1897 1088
rect 1878 1072 1881 1078
rect 2002 1068 2006 1071
rect 2018 1058 2022 1061
rect 2038 1052 2041 1108
rect 2070 1082 2073 1138
rect 2086 1092 2089 1148
rect 2114 1118 2118 1121
rect 2142 1092 2145 1168
rect 2150 1162 2153 1278
rect 2166 1242 2169 1268
rect 2198 1222 2201 1250
rect 2206 1211 2209 1328
rect 2198 1208 2209 1211
rect 2198 1132 2201 1208
rect 2214 1152 2217 1398
rect 2222 1352 2225 1398
rect 2234 1388 2238 1391
rect 2222 1222 2225 1348
rect 2246 1342 2249 1458
rect 2302 1452 2305 1548
rect 2314 1468 2318 1471
rect 2326 1462 2329 1538
rect 2438 1532 2441 1558
rect 2510 1552 2513 1658
rect 2518 1612 2521 1718
rect 2526 1662 2529 1848
rect 2542 1842 2545 1848
rect 2550 1802 2553 1868
rect 2606 1852 2609 1858
rect 2574 1822 2577 1848
rect 2598 1822 2601 1848
rect 2550 1752 2553 1758
rect 2538 1748 2542 1751
rect 2558 1751 2561 1818
rect 2582 1762 2585 1768
rect 2614 1762 2617 1858
rect 2638 1752 2641 1758
rect 2558 1748 2566 1751
rect 2578 1748 2582 1751
rect 2626 1748 2630 1751
rect 2546 1738 2550 1741
rect 2578 1738 2582 1741
rect 2550 1691 2553 1718
rect 2546 1688 2553 1691
rect 2558 1692 2561 1738
rect 2550 1672 2553 1678
rect 2574 1672 2577 1728
rect 2598 1702 2601 1748
rect 2598 1682 2601 1698
rect 2594 1678 2598 1681
rect 2542 1622 2545 1668
rect 2566 1652 2569 1668
rect 2574 1662 2577 1668
rect 2582 1662 2585 1668
rect 2506 1548 2510 1551
rect 2454 1542 2457 1548
rect 2526 1532 2529 1548
rect 2542 1532 2545 1618
rect 2586 1558 2590 1561
rect 2550 1542 2553 1548
rect 2598 1542 2601 1668
rect 2606 1622 2609 1738
rect 2638 1732 2641 1738
rect 2646 1732 2649 1768
rect 2678 1762 2681 1798
rect 2698 1768 2702 1771
rect 2710 1768 2718 1771
rect 2710 1762 2713 1768
rect 2726 1762 2729 1898
rect 2742 1892 2745 1998
rect 2830 1992 2833 2018
rect 2858 1988 2862 1991
rect 2790 1962 2793 1968
rect 2754 1958 2777 1961
rect 2774 1952 2777 1958
rect 2866 1958 2870 1961
rect 2762 1948 2766 1951
rect 2758 1872 2761 1938
rect 2766 1932 2769 1938
rect 2782 1922 2785 1928
rect 2782 1872 2785 1898
rect 2790 1892 2793 1958
rect 2814 1952 2817 1958
rect 2878 1952 2881 2008
rect 2894 1952 2897 1958
rect 2926 1952 2929 1958
rect 2858 1948 2862 1951
rect 2886 1942 2889 1948
rect 2802 1938 2806 1941
rect 2850 1938 2854 1941
rect 2934 1941 2937 2048
rect 2942 1992 2945 2058
rect 2954 1958 2958 1961
rect 2946 1948 2950 1951
rect 2934 1938 2945 1941
rect 2954 1938 2958 1941
rect 2802 1928 2806 1931
rect 2662 1742 2665 1758
rect 2678 1752 2681 1758
rect 2750 1752 2753 1848
rect 2670 1742 2673 1748
rect 2694 1742 2697 1748
rect 2726 1742 2729 1748
rect 2742 1742 2745 1748
rect 2706 1738 2710 1741
rect 2606 1542 2609 1618
rect 2614 1552 2617 1718
rect 2654 1682 2657 1698
rect 2650 1678 2654 1681
rect 2662 1672 2665 1738
rect 2670 1672 2673 1708
rect 2678 1682 2681 1688
rect 2634 1668 2638 1671
rect 2626 1658 2630 1661
rect 2642 1658 2646 1661
rect 2686 1652 2689 1708
rect 2710 1702 2713 1718
rect 2702 1662 2705 1698
rect 2622 1562 2625 1568
rect 2570 1538 2574 1541
rect 2610 1538 2617 1541
rect 2350 1472 2353 1508
rect 2366 1492 2369 1498
rect 2390 1472 2393 1498
rect 2338 1468 2342 1471
rect 2442 1468 2446 1471
rect 2294 1422 2297 1448
rect 2318 1402 2321 1458
rect 2254 1352 2257 1398
rect 2290 1368 2294 1371
rect 2326 1362 2329 1458
rect 2366 1452 2369 1468
rect 2398 1452 2401 1458
rect 2358 1432 2361 1438
rect 2358 1392 2361 1408
rect 2384 1403 2386 1407
rect 2390 1403 2393 1407
rect 2397 1403 2400 1407
rect 2358 1362 2361 1388
rect 2290 1358 2294 1361
rect 2246 1332 2249 1338
rect 2238 1271 2241 1328
rect 2254 1322 2257 1348
rect 2270 1342 2273 1358
rect 2350 1342 2353 1348
rect 2282 1338 2286 1341
rect 2322 1338 2326 1341
rect 2294 1292 2297 1318
rect 2258 1288 2262 1291
rect 2234 1268 2241 1271
rect 2238 1212 2241 1258
rect 2214 1132 2217 1138
rect 2246 1132 2249 1268
rect 2286 1262 2289 1288
rect 2270 1252 2273 1258
rect 2294 1212 2297 1268
rect 2302 1252 2305 1298
rect 2318 1262 2321 1318
rect 2326 1272 2329 1328
rect 2334 1272 2337 1298
rect 2358 1292 2361 1338
rect 2374 1312 2377 1348
rect 2382 1342 2385 1368
rect 2398 1322 2401 1348
rect 2406 1332 2409 1338
rect 2402 1318 2409 1321
rect 2374 1292 2377 1308
rect 2398 1282 2401 1308
rect 2354 1278 2377 1281
rect 2374 1272 2377 1278
rect 2362 1268 2366 1271
rect 2054 1062 2057 1078
rect 2066 1068 2070 1071
rect 2086 1062 2089 1068
rect 2094 1062 2097 1078
rect 1846 1022 1849 1050
rect 2018 1048 2022 1051
rect 2074 1048 2078 1051
rect 1854 952 1857 998
rect 1826 948 1830 951
rect 1882 948 1886 951
rect 1894 942 1897 1048
rect 2030 1042 2033 1048
rect 2102 1042 2105 1048
rect 2058 1018 2062 1021
rect 1974 1002 1977 1018
rect 1910 952 1913 968
rect 1926 952 1929 958
rect 1958 952 1961 958
rect 1982 952 1985 998
rect 2022 960 2025 979
rect 2110 952 2113 1088
rect 2158 1082 2161 1118
rect 2118 962 2121 1068
rect 2126 1032 2129 1038
rect 2134 1022 2137 1078
rect 2150 1062 2153 1078
rect 2150 992 2153 1018
rect 2158 1002 2161 1078
rect 2174 1072 2177 1078
rect 2190 1072 2193 1078
rect 2178 1058 2182 1061
rect 2150 962 2153 988
rect 1950 942 1953 948
rect 2054 942 2057 948
rect 1762 938 1766 941
rect 1850 938 1854 941
rect 1734 932 1737 938
rect 1686 808 1697 811
rect 1686 772 1689 778
rect 1634 748 1638 751
rect 1682 748 1686 751
rect 1670 742 1673 748
rect 1634 728 1638 731
rect 1670 702 1673 738
rect 1566 662 1569 668
rect 1506 648 1510 651
rect 1454 628 1465 631
rect 1430 562 1433 618
rect 1438 562 1441 598
rect 1414 542 1417 548
rect 1454 542 1457 628
rect 1462 542 1465 618
rect 1486 592 1489 618
rect 1486 552 1489 578
rect 1502 562 1505 598
rect 1534 552 1537 658
rect 1574 652 1577 678
rect 1602 668 1606 671
rect 1610 658 1614 661
rect 1590 622 1593 658
rect 1574 592 1577 608
rect 1590 592 1593 618
rect 1510 542 1513 548
rect 1542 542 1545 548
rect 1558 542 1561 558
rect 1566 552 1569 558
rect 1594 548 1598 551
rect 1474 538 1478 541
rect 1454 532 1457 538
rect 1462 532 1465 538
rect 1550 532 1553 538
rect 1434 528 1438 531
rect 1474 528 1478 531
rect 1506 528 1510 531
rect 1582 522 1585 538
rect 1438 481 1441 518
rect 1446 492 1449 508
rect 1430 478 1441 481
rect 1430 472 1433 478
rect 1418 468 1422 471
rect 1438 462 1441 468
rect 1426 458 1430 461
rect 1414 442 1417 448
rect 1446 382 1449 428
rect 1454 392 1457 468
rect 1462 462 1465 488
rect 1486 462 1489 488
rect 1518 472 1521 498
rect 1590 482 1593 548
rect 1606 541 1609 568
rect 1602 538 1609 541
rect 1614 542 1617 628
rect 1622 602 1625 678
rect 1630 642 1633 668
rect 1638 652 1641 658
rect 1658 648 1662 651
rect 1622 542 1625 548
rect 1630 542 1633 638
rect 1678 622 1681 648
rect 1654 562 1657 598
rect 1642 558 1646 561
rect 1642 538 1646 541
rect 1614 531 1617 538
rect 1614 528 1622 531
rect 1602 518 1606 521
rect 1606 482 1609 488
rect 1506 448 1510 451
rect 1474 438 1478 441
rect 1474 418 1478 421
rect 1446 352 1449 378
rect 1462 362 1465 398
rect 1398 342 1401 348
rect 1382 338 1390 341
rect 1302 322 1305 328
rect 1326 322 1329 338
rect 1378 328 1382 331
rect 1334 312 1337 318
rect 1254 262 1257 288
rect 1174 242 1177 248
rect 1182 242 1185 248
rect 1198 242 1201 248
rect 1134 162 1137 168
rect 1066 148 1073 151
rect 810 128 814 131
rect 848 103 850 107
rect 854 103 857 107
rect 861 103 864 107
rect 886 102 889 128
rect 918 82 921 98
rect 902 72 905 78
rect 958 62 961 148
rect 1054 142 1057 148
rect 970 138 974 141
rect 1014 132 1017 138
rect 1078 132 1081 158
rect 1106 148 1110 151
rect 1142 142 1145 238
rect 1158 132 1161 188
rect 1214 162 1217 218
rect 1194 158 1198 161
rect 1214 152 1217 158
rect 1230 152 1233 258
rect 1254 222 1257 248
rect 1270 182 1273 298
rect 1302 272 1305 308
rect 1318 282 1321 288
rect 1358 262 1361 308
rect 1398 292 1401 338
rect 1422 332 1425 338
rect 1398 252 1401 288
rect 1360 203 1362 207
rect 1366 203 1369 207
rect 1373 203 1376 207
rect 1270 172 1273 178
rect 1186 148 1190 151
rect 1242 148 1246 151
rect 1174 142 1177 148
rect 1202 138 1206 141
rect 1218 138 1222 141
rect 1210 128 1214 131
rect 1118 82 1121 88
rect 1102 72 1105 78
rect 1158 62 1161 68
rect 1050 58 1054 61
rect 798 22 801 48
rect 854 22 857 48
rect 1054 22 1057 48
rect 678 -22 689 -19
rect 726 -18 729 8
rect 766 -18 769 8
rect 726 -22 730 -18
rect 766 -22 770 -18
rect 1022 -19 1026 -18
rect 1030 -19 1033 18
rect 1230 12 1233 18
rect 1022 -22 1033 -19
rect 1102 -18 1105 8
rect 1214 -18 1217 8
rect 1238 -18 1241 148
rect 1262 142 1265 168
rect 1278 122 1281 178
rect 1318 162 1321 188
rect 1254 62 1257 108
rect 1302 72 1305 158
rect 1318 112 1321 148
rect 1366 142 1369 148
rect 1422 142 1425 148
rect 1382 122 1385 128
rect 1318 82 1321 88
rect 1250 58 1254 61
rect 1254 22 1257 48
rect 1254 -18 1257 8
rect 1278 -18 1281 8
rect 1360 3 1362 7
rect 1366 3 1369 7
rect 1373 3 1376 7
rect 1430 -18 1433 348
rect 1446 292 1449 318
rect 1462 271 1465 358
rect 1470 352 1473 358
rect 1478 352 1481 388
rect 1486 362 1489 438
rect 1478 322 1481 348
rect 1502 342 1505 408
rect 1518 362 1521 468
rect 1590 462 1593 468
rect 1646 462 1649 528
rect 1526 362 1529 448
rect 1526 352 1529 358
rect 1510 342 1513 348
rect 1534 342 1537 438
rect 1542 422 1545 448
rect 1550 411 1553 458
rect 1542 408 1553 411
rect 1542 362 1545 408
rect 1462 268 1473 271
rect 1470 262 1473 268
rect 1494 262 1497 318
rect 1526 292 1529 318
rect 1542 312 1545 358
rect 1550 352 1553 358
rect 1558 342 1561 448
rect 1574 352 1577 358
rect 1598 342 1601 418
rect 1606 352 1609 408
rect 1622 332 1625 398
rect 1654 382 1657 518
rect 1670 482 1673 548
rect 1686 542 1689 698
rect 1694 642 1697 808
rect 1702 762 1705 918
rect 1714 878 1718 881
rect 1710 862 1713 868
rect 1734 862 1737 908
rect 1782 892 1785 938
rect 1806 932 1809 938
rect 1798 882 1801 928
rect 1770 878 1774 881
rect 1742 872 1745 878
rect 1778 868 1782 871
rect 1778 858 1782 861
rect 1750 852 1753 858
rect 1786 848 1790 851
rect 1802 848 1806 851
rect 1718 802 1721 848
rect 1710 732 1713 798
rect 1726 752 1729 848
rect 1814 842 1817 928
rect 1830 912 1833 938
rect 1838 932 1841 938
rect 1830 862 1833 898
rect 1838 862 1841 888
rect 1846 872 1849 938
rect 1862 932 1865 938
rect 1950 932 1953 938
rect 1974 932 1977 938
rect 1870 902 1873 918
rect 1880 903 1882 907
rect 1886 903 1889 907
rect 1893 903 1896 907
rect 1918 892 1921 908
rect 1926 892 1929 918
rect 1866 888 1870 891
rect 1902 882 1905 888
rect 1942 872 1945 918
rect 1966 902 1969 928
rect 2070 912 2073 928
rect 1962 888 1966 891
rect 1734 752 1737 768
rect 1742 732 1745 738
rect 1750 732 1753 808
rect 1782 792 1785 828
rect 1814 812 1817 818
rect 1830 771 1833 858
rect 1862 802 1865 868
rect 1870 862 1873 868
rect 1882 848 1886 851
rect 1902 842 1905 868
rect 1914 858 1918 861
rect 1846 792 1849 798
rect 1830 768 1841 771
rect 1798 752 1801 758
rect 1830 752 1833 758
rect 1762 748 1766 751
rect 1806 742 1809 748
rect 1774 722 1777 738
rect 1754 718 1758 721
rect 1718 702 1721 718
rect 1742 682 1745 688
rect 1726 672 1729 678
rect 1694 592 1697 598
rect 1782 592 1785 658
rect 1826 618 1830 621
rect 1750 552 1753 588
rect 1838 562 1841 768
rect 1862 752 1865 778
rect 1894 772 1897 818
rect 1934 812 1937 848
rect 1942 842 1945 858
rect 1950 842 1953 868
rect 1998 852 2001 858
rect 2038 852 2041 878
rect 2110 872 2113 948
rect 2118 912 2121 958
rect 2166 952 2169 978
rect 2174 952 2177 1018
rect 2190 991 2193 1068
rect 2198 1062 2201 1078
rect 2198 1002 2201 1058
rect 2182 988 2193 991
rect 2174 912 2177 938
rect 2182 922 2185 988
rect 2194 978 2198 981
rect 2190 942 2193 958
rect 2202 948 2206 951
rect 2206 932 2209 938
rect 2214 882 2217 1118
rect 2254 1072 2257 1178
rect 2262 1162 2265 1188
rect 2294 1172 2297 1208
rect 2302 1192 2305 1238
rect 2310 1222 2313 1238
rect 2318 1162 2321 1218
rect 2326 1172 2329 1268
rect 2382 1262 2385 1268
rect 2398 1252 2401 1278
rect 2290 1158 2294 1161
rect 2342 1152 2345 1218
rect 2384 1203 2386 1207
rect 2390 1203 2393 1207
rect 2397 1203 2400 1207
rect 2354 1158 2358 1161
rect 2366 1152 2369 1158
rect 2306 1148 2310 1151
rect 2362 1148 2366 1151
rect 2318 1142 2321 1148
rect 2386 1138 2390 1141
rect 2310 1122 2313 1138
rect 2326 1132 2329 1138
rect 2374 1132 2377 1138
rect 2338 1118 2342 1121
rect 2234 1068 2238 1071
rect 2222 1062 2225 1068
rect 2262 1062 2265 1108
rect 2286 1082 2289 1098
rect 2302 1082 2305 1088
rect 2326 1082 2329 1088
rect 2342 1072 2345 1088
rect 2270 1062 2273 1068
rect 2230 1032 2233 1058
rect 2222 962 2225 978
rect 2230 972 2233 1028
rect 2246 962 2249 1058
rect 2262 1052 2265 1058
rect 2310 1052 2313 1068
rect 2350 1062 2353 1078
rect 2358 1072 2361 1128
rect 2362 1068 2366 1071
rect 2294 972 2297 978
rect 2342 962 2345 978
rect 2274 958 2278 961
rect 2338 958 2342 961
rect 2262 942 2265 948
rect 2278 942 2281 948
rect 2286 942 2289 958
rect 2302 942 2305 958
rect 2358 951 2361 1058
rect 2366 1042 2369 1048
rect 2382 1021 2385 1138
rect 2398 1132 2401 1138
rect 2406 1082 2409 1318
rect 2414 1262 2417 1368
rect 2430 1362 2433 1418
rect 2426 1358 2430 1361
rect 2438 1352 2441 1468
rect 2446 1442 2449 1448
rect 2438 1302 2441 1318
rect 2454 1302 2457 1528
rect 2526 1492 2529 1498
rect 2582 1482 2585 1488
rect 2606 1482 2609 1488
rect 2614 1482 2617 1538
rect 2462 1462 2465 1478
rect 2590 1472 2593 1478
rect 2474 1468 2489 1471
rect 2470 1362 2473 1458
rect 2478 1452 2481 1458
rect 2462 1342 2465 1348
rect 2478 1322 2481 1448
rect 2486 1432 2489 1468
rect 2602 1468 2606 1471
rect 2494 1452 2497 1468
rect 2510 1462 2513 1468
rect 2494 1442 2497 1448
rect 2518 1441 2521 1468
rect 2566 1462 2569 1468
rect 2542 1442 2545 1448
rect 2510 1438 2521 1441
rect 2498 1358 2502 1361
rect 2510 1342 2513 1438
rect 2534 1362 2537 1438
rect 2558 1432 2561 1458
rect 2550 1352 2553 1408
rect 2558 1402 2561 1428
rect 2566 1362 2569 1368
rect 2586 1348 2590 1351
rect 2426 1268 2430 1271
rect 2446 1262 2449 1268
rect 2462 1262 2465 1318
rect 2494 1312 2497 1338
rect 2518 1332 2521 1348
rect 2526 1342 2529 1348
rect 2558 1342 2561 1348
rect 2578 1338 2582 1341
rect 2542 1332 2545 1338
rect 2478 1292 2481 1308
rect 2534 1292 2537 1318
rect 2558 1292 2561 1338
rect 2570 1328 2574 1331
rect 2546 1278 2550 1281
rect 2486 1262 2489 1268
rect 2422 1242 2425 1258
rect 2414 1152 2417 1208
rect 2454 1192 2457 1208
rect 2462 1172 2465 1258
rect 2478 1161 2481 1218
rect 2494 1212 2497 1278
rect 2522 1258 2526 1261
rect 2510 1212 2513 1258
rect 2494 1162 2497 1168
rect 2478 1158 2489 1161
rect 2506 1158 2510 1161
rect 2442 1148 2446 1151
rect 2414 1082 2417 1148
rect 2462 1142 2465 1148
rect 2470 1142 2473 1158
rect 2478 1132 2481 1148
rect 2426 1128 2430 1131
rect 2454 1122 2457 1128
rect 2470 1118 2478 1121
rect 2454 1092 2457 1118
rect 2470 1092 2473 1118
rect 2442 1088 2446 1091
rect 2486 1071 2489 1158
rect 2518 1152 2521 1188
rect 2510 1132 2513 1138
rect 2494 1122 2497 1128
rect 2526 1122 2529 1138
rect 2498 1078 2502 1081
rect 2478 1068 2494 1071
rect 2422 1062 2425 1068
rect 2454 1062 2457 1068
rect 2374 1018 2385 1021
rect 2366 962 2369 1008
rect 2358 948 2369 951
rect 2310 942 2313 948
rect 2330 938 2334 941
rect 2222 932 2225 938
rect 2230 902 2233 938
rect 2242 918 2246 921
rect 2254 912 2257 938
rect 2262 892 2265 938
rect 2350 932 2353 948
rect 2358 932 2361 938
rect 2230 872 2233 878
rect 2294 871 2297 908
rect 2294 868 2302 871
rect 2054 862 2057 868
rect 2110 862 2113 868
rect 2174 862 2177 868
rect 2102 822 2105 848
rect 1890 768 1894 771
rect 1846 652 1849 718
rect 1880 703 1882 707
rect 1886 703 1889 707
rect 1893 703 1896 707
rect 1886 672 1889 688
rect 1858 668 1862 671
rect 1890 648 1894 651
rect 1854 642 1857 648
rect 1910 642 1913 768
rect 1934 752 1937 808
rect 2022 760 2025 779
rect 1990 742 1993 748
rect 1974 732 1977 738
rect 2054 692 2057 748
rect 2062 742 2065 818
rect 2078 762 2081 768
rect 2126 752 2129 838
rect 2134 812 2137 818
rect 2142 802 2145 858
rect 2262 831 2265 850
rect 2098 748 2102 751
rect 2130 748 2134 751
rect 2142 742 2145 798
rect 2174 752 2177 778
rect 2206 752 2209 808
rect 2214 762 2217 778
rect 2238 752 2241 798
rect 2286 781 2289 858
rect 2282 778 2289 781
rect 2294 772 2297 868
rect 2310 862 2313 888
rect 2262 752 2265 758
rect 2230 742 2233 748
rect 2082 738 2086 741
rect 2114 738 2118 741
rect 2154 738 2158 741
rect 2170 738 2174 741
rect 2290 738 2294 741
rect 2062 692 2065 738
rect 2142 728 2150 731
rect 2194 728 2198 731
rect 1962 688 1966 691
rect 1926 662 1929 668
rect 1934 652 1937 668
rect 1942 662 1945 678
rect 1950 662 1953 668
rect 1966 662 1969 678
rect 1974 672 1977 678
rect 1982 662 1985 678
rect 2046 672 2049 678
rect 2078 672 2081 728
rect 2118 701 2121 718
rect 2110 698 2121 701
rect 1994 658 1998 661
rect 1994 648 1998 651
rect 1854 562 1857 588
rect 1886 552 1889 628
rect 1910 562 1913 638
rect 1950 562 1953 638
rect 1698 548 1702 551
rect 1686 512 1689 528
rect 1686 492 1689 498
rect 1710 482 1713 538
rect 1750 532 1753 548
rect 1886 542 1889 548
rect 1914 538 1918 541
rect 1806 532 1809 538
rect 1942 532 1945 538
rect 1790 522 1793 528
rect 1750 492 1753 508
rect 1880 503 1882 507
rect 1886 503 1889 507
rect 1893 503 1896 507
rect 1782 492 1785 498
rect 1730 488 1734 491
rect 1950 491 1953 558
rect 1942 488 1953 491
rect 1974 542 1977 648
rect 2006 632 2009 668
rect 2022 662 2025 668
rect 2034 658 2038 661
rect 2054 652 2057 668
rect 2098 658 2102 661
rect 2018 648 2022 651
rect 2054 642 2057 648
rect 2014 571 2017 618
rect 2086 612 2089 648
rect 2086 592 2089 608
rect 2006 568 2025 571
rect 1974 492 1977 538
rect 1982 522 1985 558
rect 1670 422 1673 478
rect 1758 472 1761 488
rect 1786 478 1790 481
rect 1834 478 1857 481
rect 1718 452 1721 468
rect 1734 432 1737 468
rect 1782 452 1785 458
rect 1742 448 1750 451
rect 1742 432 1745 448
rect 1702 402 1705 418
rect 1638 352 1641 378
rect 1678 362 1681 388
rect 1742 372 1745 428
rect 1790 402 1793 478
rect 1814 472 1817 478
rect 1854 472 1857 478
rect 1826 468 1830 471
rect 1842 468 1846 471
rect 1838 462 1841 468
rect 1810 458 1814 461
rect 1850 458 1854 461
rect 1862 452 1865 488
rect 1918 472 1921 488
rect 1890 468 1894 471
rect 1886 462 1889 468
rect 1654 352 1657 358
rect 1686 352 1689 358
rect 1798 352 1801 418
rect 1822 392 1825 398
rect 1834 358 1838 361
rect 1726 342 1729 348
rect 1658 338 1662 341
rect 1834 338 1838 341
rect 1742 332 1745 338
rect 1586 328 1590 331
rect 1550 312 1553 318
rect 1574 292 1577 318
rect 1438 222 1441 258
rect 1462 252 1465 258
rect 1502 252 1505 278
rect 1518 272 1521 278
rect 1534 272 1537 278
rect 1510 262 1513 268
rect 1566 262 1569 288
rect 1594 268 1598 271
rect 1618 268 1622 271
rect 1582 262 1585 268
rect 1630 262 1633 288
rect 1654 262 1657 278
rect 1682 268 1686 271
rect 1542 252 1545 258
rect 1578 248 1590 251
rect 1534 242 1537 248
rect 1614 242 1617 258
rect 1626 248 1630 251
rect 1638 242 1641 248
rect 1490 238 1494 241
rect 1562 238 1566 241
rect 1634 218 1638 221
rect 1458 188 1462 191
rect 1478 182 1481 218
rect 1566 162 1569 218
rect 1522 148 1526 151
rect 1462 92 1465 128
rect 1486 72 1489 118
rect 1518 72 1521 98
rect 1526 82 1529 148
rect 1582 142 1585 218
rect 1662 192 1665 268
rect 1670 252 1673 258
rect 1686 231 1689 258
rect 1694 252 1697 328
rect 1726 262 1729 278
rect 1754 268 1758 271
rect 1702 252 1705 258
rect 1718 241 1721 248
rect 1714 238 1721 241
rect 1686 228 1697 231
rect 1630 162 1633 188
rect 1654 172 1657 178
rect 1566 102 1569 128
rect 1526 62 1529 68
rect 1566 62 1569 78
rect 1614 72 1617 88
rect 1630 72 1633 78
rect 1694 52 1697 228
rect 1702 182 1705 218
rect 1734 202 1737 268
rect 1742 252 1745 258
rect 1758 252 1761 258
rect 1766 252 1769 308
rect 1798 262 1801 278
rect 1818 268 1822 271
rect 1774 252 1777 258
rect 1790 241 1793 248
rect 1786 238 1793 241
rect 1806 232 1809 268
rect 1830 262 1833 308
rect 1846 271 1849 428
rect 1870 372 1873 378
rect 1854 362 1857 368
rect 1886 352 1889 438
rect 1894 432 1897 458
rect 1894 362 1897 368
rect 1862 342 1865 348
rect 1862 292 1865 328
rect 1870 302 1873 348
rect 1880 303 1882 307
rect 1886 303 1889 307
rect 1893 303 1896 307
rect 1902 272 1905 388
rect 1910 332 1913 448
rect 1934 441 1937 468
rect 1942 462 1945 488
rect 1950 472 1953 478
rect 1982 472 1985 478
rect 1942 452 1945 458
rect 1966 448 1974 451
rect 1934 438 1945 441
rect 1934 372 1937 408
rect 1942 392 1945 438
rect 1922 328 1926 331
rect 1934 292 1937 368
rect 1950 342 1953 398
rect 1966 392 1969 448
rect 1990 402 1993 418
rect 1998 392 2001 548
rect 2006 542 2009 568
rect 2022 562 2025 568
rect 2062 562 2065 588
rect 2110 571 2113 698
rect 2118 682 2121 688
rect 2142 672 2145 728
rect 2158 672 2161 698
rect 2174 682 2177 688
rect 2130 658 2134 661
rect 2146 658 2150 661
rect 2134 642 2137 648
rect 2102 568 2113 571
rect 2126 638 2134 641
rect 2014 552 2017 558
rect 2102 552 2105 568
rect 2126 562 2129 638
rect 2166 622 2169 668
rect 2182 662 2185 668
rect 2110 552 2113 558
rect 2134 552 2137 608
rect 2166 552 2169 558
rect 2014 452 2017 548
rect 2046 542 2049 548
rect 2082 538 2086 541
rect 2138 538 2142 541
rect 2062 532 2065 538
rect 2118 532 2121 538
rect 2074 528 2078 531
rect 2142 522 2145 538
rect 2162 528 2166 531
rect 2030 462 2033 518
rect 2054 512 2057 518
rect 2070 482 2073 488
rect 2086 472 2089 478
rect 2142 472 2145 518
rect 2030 382 2033 458
rect 2118 422 2121 450
rect 2126 402 2129 458
rect 2090 368 2094 371
rect 2030 362 2033 368
rect 2102 362 2105 378
rect 1974 342 1977 358
rect 1982 352 1985 358
rect 2006 342 2009 358
rect 2126 352 2129 398
rect 2026 348 2030 351
rect 2082 348 2086 351
rect 1926 272 1929 288
rect 1842 268 1849 271
rect 1878 262 1881 268
rect 1950 262 1953 338
rect 1990 332 1993 338
rect 1958 312 1961 328
rect 1958 272 1961 308
rect 1970 278 1974 281
rect 1990 272 1993 318
rect 1998 292 2001 318
rect 2014 272 2017 348
rect 2062 342 2065 348
rect 2026 338 2030 341
rect 2082 338 2086 341
rect 2022 328 2030 331
rect 2022 292 2025 328
rect 2030 272 2033 278
rect 2038 272 2041 328
rect 2046 312 2049 338
rect 2110 332 2113 338
rect 2058 328 2062 331
rect 2106 328 2110 331
rect 2138 328 2142 331
rect 2070 292 2073 318
rect 2150 291 2153 518
rect 2158 472 2161 478
rect 2166 462 2169 478
rect 2182 462 2185 518
rect 2190 482 2193 648
rect 2198 612 2201 698
rect 2214 612 2217 718
rect 2198 542 2201 608
rect 2206 542 2209 548
rect 2222 541 2225 708
rect 2230 662 2233 738
rect 2254 672 2257 718
rect 2302 702 2305 718
rect 2278 672 2281 688
rect 2294 672 2297 678
rect 2310 671 2313 858
rect 2318 752 2321 908
rect 2366 901 2369 948
rect 2374 912 2377 1018
rect 2430 1012 2433 1058
rect 2442 1048 2446 1051
rect 2462 1012 2465 1068
rect 2384 1003 2386 1007
rect 2390 1003 2393 1007
rect 2397 1003 2400 1007
rect 2470 982 2473 1048
rect 2382 952 2385 958
rect 2390 942 2393 968
rect 2478 962 2481 1068
rect 2518 1062 2521 1078
rect 2526 1062 2529 1068
rect 2534 1062 2537 1148
rect 2542 1132 2545 1138
rect 2550 1081 2553 1158
rect 2558 1132 2561 1278
rect 2574 1262 2577 1268
rect 2566 1252 2569 1258
rect 2590 1172 2593 1218
rect 2598 1162 2601 1468
rect 2614 1462 2617 1468
rect 2606 1392 2609 1438
rect 2622 1282 2625 1558
rect 2634 1548 2638 1551
rect 2646 1542 2649 1588
rect 2654 1562 2657 1568
rect 2662 1542 2665 1638
rect 2670 1592 2673 1648
rect 2686 1592 2689 1648
rect 2710 1622 2713 1668
rect 2718 1662 2721 1668
rect 2726 1662 2729 1678
rect 2734 1652 2737 1738
rect 2742 1732 2745 1738
rect 2758 1712 2761 1868
rect 2790 1862 2793 1868
rect 2814 1862 2817 1908
rect 2838 1882 2841 1918
rect 2846 1902 2849 1938
rect 2886 1922 2889 1938
rect 2850 1878 2854 1881
rect 2822 1872 2825 1878
rect 2774 1852 2777 1858
rect 2830 1852 2833 1858
rect 2794 1848 2798 1851
rect 2810 1848 2814 1851
rect 2766 1762 2769 1818
rect 2838 1802 2841 1878
rect 2846 1862 2849 1868
rect 2806 1762 2809 1798
rect 2770 1758 2774 1761
rect 2822 1752 2825 1798
rect 2862 1771 2865 1898
rect 2878 1872 2881 1878
rect 2894 1862 2897 1928
rect 2902 1922 2905 1928
rect 2904 1903 2906 1907
rect 2910 1903 2913 1907
rect 2917 1903 2920 1907
rect 2942 1892 2945 1938
rect 2958 1922 2961 1928
rect 2966 1922 2969 2078
rect 2986 2068 2990 2071
rect 3022 2062 3025 2108
rect 3038 2082 3041 2138
rect 3090 2128 3094 2131
rect 3046 2092 3049 2118
rect 3054 2082 3057 2128
rect 2974 2052 2977 2058
rect 3030 2052 3033 2068
rect 3006 2042 3009 2048
rect 3038 2042 3041 2078
rect 3054 2072 3057 2078
rect 3050 2058 3054 2061
rect 3062 2042 3065 2128
rect 3094 2082 3097 2088
rect 3118 2072 3121 2158
rect 3154 2148 3158 2151
rect 3126 2112 3129 2148
rect 3142 2138 3150 2141
rect 3126 2092 3129 2108
rect 3134 2102 3137 2138
rect 3134 2072 3137 2098
rect 3142 2092 3145 2138
rect 3154 2128 3158 2131
rect 3154 2078 3158 2081
rect 3166 2072 3169 2098
rect 3174 2092 3177 2268
rect 3190 2261 3193 2338
rect 3206 2331 3209 2338
rect 3202 2328 3209 2331
rect 3230 2332 3233 2338
rect 3242 2328 3246 2331
rect 3222 2302 3225 2318
rect 3230 2302 3233 2318
rect 3226 2288 3230 2291
rect 3202 2268 3206 2271
rect 3226 2268 3230 2271
rect 3182 2258 3193 2261
rect 3210 2258 3214 2261
rect 3182 2142 3185 2258
rect 3190 2162 3193 2248
rect 3222 2222 3225 2228
rect 3198 2162 3201 2178
rect 3214 2152 3217 2158
rect 3190 2131 3193 2148
rect 3222 2142 3225 2218
rect 3230 2142 3233 2148
rect 3186 2128 3193 2131
rect 3186 2078 3190 2081
rect 3114 2058 3118 2061
rect 3130 2058 3134 2061
rect 3086 2052 3089 2058
rect 2982 1962 2985 2018
rect 2982 1952 2985 1958
rect 2974 1942 2977 1948
rect 2998 1942 3001 1998
rect 3014 1992 3017 2038
rect 3022 1942 3025 1958
rect 3034 1948 3038 1951
rect 3050 1948 3057 1951
rect 3066 1948 3070 1951
rect 3054 1942 3057 1948
rect 3078 1942 3081 1948
rect 2978 1938 2985 1941
rect 2922 1878 2926 1881
rect 2950 1872 2953 1908
rect 2958 1882 2961 1918
rect 2982 1892 2985 1938
rect 3066 1938 3070 1941
rect 2990 1932 2993 1938
rect 2998 1932 3001 1938
rect 2938 1868 2942 1871
rect 2978 1868 2982 1871
rect 2874 1858 2878 1861
rect 2894 1772 2897 1858
rect 2934 1852 2937 1858
rect 2946 1848 2950 1851
rect 2986 1848 2990 1851
rect 2862 1768 2873 1771
rect 2882 1768 2886 1771
rect 2850 1758 2854 1761
rect 2862 1752 2865 1758
rect 2794 1748 2798 1751
rect 2870 1742 2873 1768
rect 2878 1742 2881 1748
rect 2778 1738 2782 1741
rect 2826 1738 2830 1741
rect 2766 1672 2769 1698
rect 2790 1692 2793 1738
rect 2870 1702 2873 1738
rect 2786 1678 2790 1681
rect 2798 1672 2801 1698
rect 2870 1682 2873 1698
rect 2886 1682 2889 1758
rect 2918 1732 2921 1758
rect 2942 1752 2945 1788
rect 2950 1762 2953 1838
rect 2938 1738 2942 1741
rect 2950 1712 2953 1758
rect 2904 1703 2906 1707
rect 2910 1703 2913 1707
rect 2917 1703 2920 1707
rect 2926 1682 2929 1688
rect 2850 1678 2854 1681
rect 2814 1672 2817 1678
rect 2866 1668 2870 1671
rect 2830 1662 2833 1668
rect 2778 1658 2782 1661
rect 2818 1658 2825 1661
rect 2822 1652 2825 1658
rect 2838 1652 2841 1668
rect 2870 1652 2873 1658
rect 2746 1648 2750 1651
rect 2734 1622 2737 1648
rect 2702 1572 2705 1618
rect 2750 1602 2753 1618
rect 2646 1522 2649 1538
rect 2630 1470 2633 1471
rect 2634 1466 2638 1469
rect 2618 1258 2622 1261
rect 2614 1232 2617 1238
rect 2622 1192 2625 1218
rect 2614 1152 2617 1168
rect 2630 1152 2633 1466
rect 2646 1451 2649 1468
rect 2638 1448 2649 1451
rect 2662 1451 2665 1538
rect 2678 1472 2681 1478
rect 2710 1472 2713 1488
rect 2678 1452 2681 1458
rect 2658 1448 2665 1451
rect 2726 1451 2729 1548
rect 2766 1532 2769 1578
rect 2814 1562 2817 1648
rect 2830 1562 2833 1588
rect 2854 1562 2857 1568
rect 2782 1532 2785 1538
rect 2734 1462 2737 1508
rect 2742 1472 2745 1498
rect 2750 1482 2753 1508
rect 2750 1472 2753 1478
rect 2758 1452 2761 1458
rect 2782 1452 2785 1518
rect 2806 1472 2809 1508
rect 2846 1502 2849 1558
rect 2870 1552 2873 1568
rect 2878 1552 2881 1608
rect 2886 1602 2889 1678
rect 2918 1672 2921 1678
rect 2910 1662 2913 1668
rect 2894 1572 2897 1578
rect 2918 1572 2921 1668
rect 2958 1662 2961 1828
rect 2982 1812 2985 1848
rect 2990 1752 2993 1838
rect 2970 1748 2974 1751
rect 2970 1738 2974 1741
rect 2974 1722 2977 1728
rect 2974 1692 2977 1708
rect 2982 1682 2985 1688
rect 2970 1668 2974 1671
rect 2982 1662 2985 1668
rect 2990 1662 2993 1748
rect 2998 1742 3001 1868
rect 3006 1812 3009 1938
rect 3038 1912 3041 1938
rect 3046 1902 3049 1918
rect 3014 1892 3017 1898
rect 3062 1892 3065 1898
rect 3046 1882 3049 1888
rect 3086 1882 3089 2038
rect 3094 1962 3097 2018
rect 3102 1942 3105 2028
rect 3110 1942 3113 1948
rect 3026 1858 3030 1861
rect 3038 1851 3041 1878
rect 3030 1848 3041 1851
rect 2998 1672 3001 1738
rect 3006 1732 3009 1738
rect 3022 1692 3025 1798
rect 3030 1762 3033 1848
rect 3054 1812 3057 1858
rect 3070 1792 3073 1848
rect 3078 1812 3081 1868
rect 3086 1842 3089 1878
rect 3094 1872 3097 1918
rect 3102 1892 3105 1918
rect 3110 1882 3113 1908
rect 3030 1742 3033 1758
rect 3082 1748 3086 1751
rect 3094 1742 3097 1748
rect 3110 1742 3113 1878
rect 3118 1862 3121 2048
rect 3158 1982 3161 2058
rect 3182 1971 3185 2078
rect 3198 2072 3201 2098
rect 3206 2092 3209 2138
rect 3214 2082 3217 2128
rect 3222 2108 3230 2111
rect 3222 2082 3225 2108
rect 3238 2082 3241 2328
rect 3262 2272 3265 2338
rect 3270 2332 3273 2478
rect 3278 2442 3281 2448
rect 3278 2342 3281 2438
rect 3286 2392 3289 2478
rect 3294 2472 3297 2478
rect 3302 2462 3305 2488
rect 3310 2482 3313 2508
rect 3294 2352 3297 2398
rect 3290 2338 3294 2341
rect 3282 2278 3286 2281
rect 3270 2272 3273 2278
rect 3302 2272 3305 2358
rect 3298 2258 3302 2261
rect 3246 2232 3249 2258
rect 3246 2162 3249 2168
rect 3254 2162 3257 2248
rect 3270 2152 3273 2168
rect 3258 2148 3262 2151
rect 3278 2151 3281 2218
rect 3298 2158 3302 2161
rect 3278 2148 3286 2151
rect 3294 2142 3297 2148
rect 3250 2138 3254 2141
rect 3246 2112 3249 2118
rect 3246 2072 3249 2078
rect 3226 2058 3230 2061
rect 3190 2022 3193 2058
rect 3238 2052 3241 2058
rect 3262 2052 3265 2058
rect 3270 2052 3273 2098
rect 3278 2092 3281 2138
rect 3302 2082 3305 2158
rect 3310 2142 3313 2408
rect 3318 2152 3321 2518
rect 3326 2462 3329 2488
rect 3334 2472 3337 2518
rect 3366 2492 3369 2538
rect 3382 2492 3385 2618
rect 3398 2562 3401 2648
rect 3406 2632 3409 2678
rect 3422 2652 3425 2658
rect 3408 2603 3410 2607
rect 3414 2603 3417 2607
rect 3421 2603 3424 2607
rect 3438 2572 3441 2618
rect 3398 2552 3401 2558
rect 3446 2552 3449 2658
rect 3454 2622 3457 2678
rect 3474 2668 3486 2671
rect 3470 2652 3473 2658
rect 3470 2562 3473 2648
rect 3478 2552 3481 2568
rect 3494 2562 3497 2648
rect 3502 2632 3505 2738
rect 3590 2732 3593 2748
rect 3614 2738 3622 2741
rect 3530 2728 3534 2731
rect 3526 2672 3529 2718
rect 3542 2712 3545 2718
rect 3582 2702 3585 2718
rect 3542 2662 3545 2698
rect 3566 2662 3569 2688
rect 3590 2682 3593 2688
rect 3514 2648 3518 2651
rect 3562 2648 3566 2651
rect 3534 2642 3537 2648
rect 3574 2642 3577 2658
rect 3590 2642 3593 2648
rect 3566 2632 3569 2638
rect 3502 2612 3505 2618
rect 3526 2592 3529 2618
rect 3494 2552 3497 2558
rect 3518 2552 3521 2558
rect 3446 2542 3449 2548
rect 3494 2532 3497 2548
rect 3502 2542 3505 2548
rect 3526 2542 3529 2578
rect 3598 2572 3601 2718
rect 3614 2672 3617 2718
rect 3630 2692 3633 2748
rect 3630 2672 3633 2678
rect 3638 2672 3641 2718
rect 3606 2662 3609 2668
rect 3630 2662 3633 2668
rect 3626 2648 3630 2651
rect 3646 2621 3649 2738
rect 3654 2682 3657 2758
rect 3662 2742 3665 2758
rect 3706 2748 3710 2751
rect 3670 2742 3673 2748
rect 3742 2732 3745 2738
rect 3750 2732 3753 2758
rect 3758 2742 3761 2748
rect 3774 2742 3777 2808
rect 3774 2732 3777 2738
rect 3750 2722 3753 2728
rect 3682 2718 3686 2721
rect 3670 2682 3673 2698
rect 3710 2682 3713 2708
rect 3698 2678 3702 2681
rect 3658 2658 3662 2661
rect 3706 2658 3710 2661
rect 3730 2658 3734 2661
rect 3658 2648 3662 2651
rect 3638 2618 3649 2621
rect 3590 2562 3593 2568
rect 3614 2562 3617 2568
rect 3546 2558 3550 2561
rect 3542 2542 3545 2548
rect 3402 2528 3406 2531
rect 3458 2528 3462 2531
rect 3574 2522 3577 2548
rect 3398 2512 3401 2518
rect 3394 2478 3398 2481
rect 3366 2472 3369 2478
rect 3414 2472 3417 2518
rect 3386 2468 3390 2471
rect 3402 2468 3406 2471
rect 3374 2462 3377 2468
rect 3342 2452 3345 2458
rect 3326 2352 3329 2438
rect 3326 2242 3329 2348
rect 3334 2332 3337 2448
rect 3350 2372 3353 2458
rect 3362 2448 3366 2451
rect 3394 2448 3398 2451
rect 3414 2432 3417 2458
rect 3342 2352 3345 2358
rect 3358 2351 3361 2428
rect 3354 2348 3361 2351
rect 3342 2282 3345 2318
rect 3334 2262 3337 2268
rect 3326 2152 3329 2228
rect 3334 2192 3337 2258
rect 3350 2251 3353 2348
rect 3358 2332 3361 2338
rect 3366 2282 3369 2418
rect 3408 2403 3410 2407
rect 3414 2403 3417 2407
rect 3421 2403 3424 2407
rect 3438 2372 3441 2488
rect 3446 2462 3449 2468
rect 3466 2448 3470 2451
rect 3478 2442 3481 2508
rect 3494 2472 3497 2518
rect 3518 2482 3521 2518
rect 3542 2491 3545 2518
rect 3542 2488 3553 2491
rect 3486 2462 3489 2468
rect 3518 2462 3521 2468
rect 3498 2448 3502 2451
rect 3530 2448 3534 2451
rect 3542 2442 3545 2478
rect 3550 2462 3553 2488
rect 3562 2478 3566 2481
rect 3586 2478 3590 2481
rect 3606 2462 3609 2558
rect 3638 2552 3641 2618
rect 3646 2562 3649 2578
rect 3670 2552 3673 2598
rect 3614 2542 3617 2548
rect 3662 2542 3665 2548
rect 3678 2542 3681 2618
rect 3710 2592 3713 2648
rect 3694 2562 3697 2568
rect 3686 2552 3689 2558
rect 3642 2538 3646 2541
rect 3614 2462 3617 2468
rect 3578 2458 3582 2461
rect 3446 2432 3449 2438
rect 3510 2432 3513 2438
rect 3550 2431 3553 2448
rect 3542 2428 3553 2431
rect 3622 2432 3625 2538
rect 3630 2492 3633 2508
rect 3654 2502 3657 2518
rect 3670 2512 3673 2538
rect 3702 2532 3705 2578
rect 3726 2552 3729 2628
rect 3734 2561 3737 2618
rect 3758 2562 3761 2568
rect 3774 2562 3777 2648
rect 3734 2558 3742 2561
rect 3762 2548 3766 2551
rect 3746 2538 3750 2541
rect 3718 2512 3721 2538
rect 3386 2348 3390 2351
rect 3362 2268 3366 2271
rect 3374 2261 3377 2348
rect 3406 2332 3409 2358
rect 3446 2352 3449 2368
rect 3462 2362 3465 2368
rect 3454 2342 3457 2358
rect 3470 2352 3473 2418
rect 3418 2318 3422 2321
rect 3486 2282 3489 2318
rect 3434 2278 3438 2281
rect 3458 2278 3462 2281
rect 3458 2268 3462 2271
rect 3482 2268 3486 2271
rect 3398 2262 3401 2268
rect 3374 2258 3382 2261
rect 3386 2258 3390 2261
rect 3358 2252 3361 2258
rect 3350 2248 3358 2251
rect 3430 2242 3433 2248
rect 3374 2152 3377 2238
rect 3398 2182 3401 2218
rect 3408 2203 3410 2207
rect 3414 2203 3417 2207
rect 3421 2203 3424 2207
rect 3390 2162 3393 2168
rect 3406 2152 3409 2188
rect 3430 2162 3433 2238
rect 3454 2192 3457 2258
rect 3478 2252 3481 2258
rect 3486 2241 3489 2258
rect 3482 2238 3489 2241
rect 3494 2222 3497 2328
rect 3510 2262 3513 2348
rect 3518 2302 3521 2418
rect 3526 2352 3529 2388
rect 3542 2362 3545 2428
rect 3550 2392 3553 2418
rect 3542 2332 3545 2358
rect 3550 2332 3553 2378
rect 3582 2352 3585 2418
rect 3598 2362 3601 2368
rect 3598 2352 3601 2358
rect 3562 2348 3566 2351
rect 3594 2338 3598 2341
rect 3606 2332 3609 2418
rect 3622 2392 3625 2398
rect 3614 2372 3617 2378
rect 3630 2362 3633 2448
rect 3614 2342 3617 2348
rect 3630 2342 3633 2358
rect 3622 2338 3630 2341
rect 3542 2312 3545 2318
rect 3570 2288 3574 2291
rect 3518 2282 3521 2288
rect 3574 2272 3577 2278
rect 3526 2262 3529 2268
rect 3534 2262 3537 2268
rect 3510 2242 3513 2248
rect 3518 2232 3521 2258
rect 3534 2252 3537 2258
rect 3510 2192 3513 2218
rect 3542 2192 3545 2268
rect 3582 2262 3585 2308
rect 3550 2252 3553 2258
rect 3590 2252 3593 2308
rect 3610 2258 3614 2261
rect 3622 2252 3625 2338
rect 3638 2332 3641 2498
rect 3734 2492 3737 2538
rect 3774 2512 3777 2558
rect 3694 2472 3697 2478
rect 3702 2472 3705 2478
rect 3750 2472 3753 2478
rect 3646 2462 3649 2468
rect 3694 2442 3697 2468
rect 3702 2462 3705 2468
rect 3674 2418 3678 2421
rect 3662 2372 3665 2388
rect 3670 2382 3673 2388
rect 3702 2372 3705 2378
rect 3734 2372 3737 2418
rect 3742 2372 3745 2398
rect 3686 2352 3689 2358
rect 3710 2352 3713 2368
rect 3746 2358 3750 2361
rect 3562 2248 3566 2251
rect 3314 2128 3318 2131
rect 3334 2102 3337 2138
rect 3342 2132 3345 2148
rect 3342 2082 3345 2108
rect 3294 2072 3297 2078
rect 3182 1968 3193 1971
rect 3178 1958 3182 1961
rect 3150 1952 3153 1958
rect 3150 1942 3153 1948
rect 3158 1942 3161 1948
rect 3170 1938 3174 1941
rect 3138 1928 3142 1931
rect 3126 1912 3129 1918
rect 3118 1832 3121 1858
rect 3134 1842 3137 1888
rect 3150 1872 3153 1938
rect 3190 1932 3193 1968
rect 3214 1952 3217 2008
rect 3262 1992 3265 2018
rect 3158 1872 3161 1898
rect 3142 1862 3145 1868
rect 3166 1862 3169 1868
rect 3182 1862 3185 1918
rect 3198 1872 3201 1918
rect 3206 1912 3209 1938
rect 3222 1932 3225 1988
rect 3238 1952 3241 1958
rect 3262 1952 3265 1958
rect 3274 1948 3278 1951
rect 3278 1932 3281 1938
rect 3286 1932 3289 2008
rect 3294 1972 3297 2068
rect 3302 2062 3305 2068
rect 3318 2062 3321 2068
rect 3310 2052 3313 2058
rect 3334 2052 3337 2078
rect 3310 2022 3313 2048
rect 3302 2018 3310 2021
rect 3302 1952 3305 2018
rect 3310 1952 3313 1958
rect 3326 1952 3329 2018
rect 3338 1948 3342 1951
rect 3302 1932 3305 1938
rect 3222 1901 3225 1928
rect 3218 1898 3225 1901
rect 3210 1888 3214 1891
rect 3154 1848 3158 1851
rect 3170 1848 3174 1851
rect 3186 1848 3190 1851
rect 3214 1842 3217 1868
rect 3230 1862 3233 1898
rect 3238 1882 3241 1908
rect 3246 1892 3249 1918
rect 3254 1912 3257 1928
rect 3254 1882 3257 1898
rect 3286 1882 3289 1898
rect 3310 1882 3313 1938
rect 3330 1928 3334 1931
rect 3318 1882 3321 1928
rect 3334 1882 3337 1908
rect 3242 1878 3246 1881
rect 3302 1872 3305 1878
rect 3334 1872 3337 1878
rect 3274 1868 3278 1871
rect 3242 1858 3246 1861
rect 3274 1858 3278 1861
rect 3306 1858 3310 1861
rect 3338 1858 3342 1861
rect 3118 1752 3121 1768
rect 3126 1752 3129 1818
rect 3198 1792 3201 1838
rect 3222 1832 3225 1858
rect 3258 1848 3262 1851
rect 3166 1772 3169 1778
rect 3134 1752 3137 1758
rect 3114 1738 3121 1741
rect 3010 1678 3014 1681
rect 3030 1662 3033 1738
rect 3082 1728 3089 1731
rect 3058 1718 3062 1721
rect 3046 1692 3049 1718
rect 3078 1692 3081 1708
rect 2942 1582 2945 1648
rect 2990 1612 2993 1658
rect 2942 1562 2945 1578
rect 2886 1542 2889 1558
rect 2910 1552 2913 1558
rect 2874 1538 2878 1541
rect 2854 1522 2857 1528
rect 2814 1482 2817 1488
rect 2838 1472 2841 1488
rect 2846 1472 2849 1498
rect 2854 1462 2857 1498
rect 2886 1492 2889 1508
rect 2798 1452 2801 1458
rect 2726 1448 2737 1451
rect 2846 1451 2849 1458
rect 2846 1448 2854 1451
rect 2638 1252 2641 1448
rect 2654 1442 2657 1448
rect 2670 1442 2673 1448
rect 2686 1442 2689 1448
rect 2718 1432 2721 1448
rect 2646 1322 2649 1348
rect 2702 1342 2705 1418
rect 2734 1352 2737 1448
rect 2774 1421 2777 1448
rect 2814 1441 2817 1448
rect 2802 1438 2817 1441
rect 2870 1422 2873 1448
rect 2894 1422 2897 1548
rect 2934 1542 2937 1548
rect 2966 1532 2969 1558
rect 2982 1542 2985 1568
rect 2998 1562 3001 1578
rect 2994 1548 2998 1551
rect 2974 1522 2977 1528
rect 2904 1503 2906 1507
rect 2910 1503 2913 1507
rect 2917 1503 2920 1507
rect 2942 1462 2945 1468
rect 2774 1418 2785 1421
rect 2750 1362 2753 1388
rect 2758 1362 2761 1418
rect 2770 1358 2774 1361
rect 2686 1322 2689 1328
rect 2646 1292 2649 1298
rect 2686 1262 2689 1308
rect 2726 1282 2729 1288
rect 2742 1272 2745 1278
rect 2774 1272 2777 1318
rect 2782 1302 2785 1418
rect 2846 1412 2849 1418
rect 2790 1352 2793 1368
rect 2802 1358 2806 1361
rect 2846 1361 2849 1408
rect 2854 1372 2857 1378
rect 2842 1358 2849 1361
rect 2810 1348 2814 1351
rect 2838 1342 2841 1348
rect 2822 1338 2830 1341
rect 2798 1312 2801 1338
rect 2814 1272 2817 1298
rect 2822 1292 2825 1338
rect 2838 1322 2841 1338
rect 2826 1288 2830 1291
rect 2830 1272 2833 1278
rect 2642 1248 2646 1251
rect 2646 1192 2649 1198
rect 2686 1152 2689 1258
rect 2774 1222 2777 1250
rect 2790 1162 2793 1188
rect 2742 1142 2745 1158
rect 2822 1152 2825 1168
rect 2574 1132 2577 1138
rect 2566 1121 2569 1128
rect 2566 1118 2582 1121
rect 2542 1078 2553 1081
rect 2558 1082 2561 1088
rect 2542 1072 2545 1078
rect 2582 1072 2585 1108
rect 2590 1092 2593 1118
rect 2598 1112 2601 1128
rect 2606 1112 2609 1128
rect 2638 1122 2641 1128
rect 2598 1082 2601 1088
rect 2606 1072 2609 1078
rect 2542 1062 2545 1068
rect 2490 1058 2494 1061
rect 2494 952 2497 968
rect 2502 952 2505 1048
rect 2418 948 2422 951
rect 2474 948 2478 951
rect 2502 942 2505 948
rect 2510 942 2513 1018
rect 2526 952 2529 958
rect 2538 948 2542 951
rect 2442 938 2446 941
rect 2450 928 2454 931
rect 2366 898 2377 901
rect 2338 878 2342 881
rect 2358 872 2361 898
rect 2374 892 2377 898
rect 2366 872 2369 878
rect 2342 858 2350 861
rect 2326 822 2329 848
rect 2326 802 2329 818
rect 2342 792 2345 858
rect 2390 852 2393 928
rect 2462 921 2465 938
rect 2478 932 2481 938
rect 2454 918 2465 921
rect 2402 888 2406 891
rect 2430 882 2433 918
rect 2446 892 2449 898
rect 2438 882 2441 888
rect 2454 872 2457 918
rect 2486 902 2489 938
rect 2534 932 2537 938
rect 2382 842 2385 848
rect 2366 792 2369 828
rect 2384 803 2386 807
rect 2390 803 2393 807
rect 2397 803 2400 807
rect 2318 692 2321 748
rect 2326 742 2329 748
rect 2334 742 2337 768
rect 2358 762 2361 778
rect 2342 731 2345 748
rect 2334 728 2345 731
rect 2302 668 2313 671
rect 2334 672 2337 728
rect 2350 672 2353 678
rect 2262 662 2265 668
rect 2286 662 2289 668
rect 2302 662 2305 668
rect 2358 662 2361 758
rect 2374 732 2377 798
rect 2414 742 2417 858
rect 2422 832 2425 858
rect 2430 852 2433 868
rect 2454 862 2457 868
rect 2462 862 2465 898
rect 2510 882 2513 928
rect 2518 912 2521 918
rect 2474 878 2478 881
rect 2522 878 2526 881
rect 2486 872 2489 878
rect 2494 862 2497 868
rect 2462 852 2465 858
rect 2510 842 2513 878
rect 2534 862 2537 898
rect 2550 892 2553 1068
rect 2578 1058 2582 1061
rect 2566 1052 2569 1058
rect 2558 962 2561 968
rect 2566 962 2569 968
rect 2582 952 2585 958
rect 2590 952 2593 1038
rect 2598 972 2601 1068
rect 2606 1052 2609 1068
rect 2630 1062 2633 1118
rect 2650 1088 2654 1091
rect 2638 1072 2641 1078
rect 2662 1062 2665 1128
rect 2726 1122 2729 1128
rect 2678 1072 2681 1088
rect 2710 1072 2713 1078
rect 2742 1072 2745 1098
rect 2758 1082 2761 1088
rect 2618 1058 2622 1061
rect 2630 952 2633 1058
rect 2646 1052 2649 1058
rect 2670 982 2673 1068
rect 2686 1062 2689 1068
rect 2718 1062 2721 1068
rect 2734 1052 2737 1058
rect 2698 1048 2702 1051
rect 2706 1048 2713 1051
rect 2722 1048 2726 1051
rect 2670 972 2673 978
rect 2642 958 2646 961
rect 2654 952 2657 958
rect 2686 952 2689 1018
rect 2626 948 2630 951
rect 2578 938 2582 941
rect 2602 938 2606 941
rect 2666 938 2670 941
rect 2558 912 2561 918
rect 2590 912 2593 938
rect 2646 932 2649 938
rect 2686 932 2689 938
rect 2618 928 2622 931
rect 2542 842 2545 878
rect 2558 862 2561 898
rect 2430 762 2433 768
rect 2422 742 2425 748
rect 2410 738 2414 741
rect 2402 728 2406 731
rect 2366 682 2369 718
rect 2406 671 2409 718
rect 2402 668 2409 671
rect 2430 672 2433 758
rect 2454 752 2457 768
rect 2438 732 2441 738
rect 2446 702 2449 748
rect 2454 732 2457 738
rect 2450 688 2454 691
rect 2438 662 2441 688
rect 2462 672 2465 808
rect 2478 742 2481 818
rect 2494 792 2497 828
rect 2518 762 2521 788
rect 2526 782 2529 818
rect 2550 802 2553 818
rect 2566 812 2569 878
rect 2606 872 2609 878
rect 2614 872 2617 918
rect 2638 872 2641 878
rect 2662 872 2665 918
rect 2702 882 2705 918
rect 2682 878 2686 881
rect 2586 868 2590 871
rect 2690 868 2694 871
rect 2622 862 2625 868
rect 2630 862 2633 868
rect 2670 862 2673 868
rect 2682 858 2686 861
rect 2582 772 2585 858
rect 2614 812 2617 858
rect 2490 748 2494 751
rect 2514 748 2518 751
rect 2490 738 2494 741
rect 2474 728 2478 731
rect 2486 692 2489 728
rect 2338 658 2342 661
rect 2238 602 2241 618
rect 2234 558 2238 561
rect 2246 552 2249 658
rect 2254 622 2257 658
rect 2302 652 2305 658
rect 2310 652 2313 658
rect 2354 648 2358 651
rect 2282 618 2286 621
rect 2318 612 2321 648
rect 2270 572 2273 608
rect 2326 602 2329 648
rect 2266 568 2270 571
rect 2242 548 2246 551
rect 2222 538 2230 541
rect 2214 532 2217 538
rect 2166 342 2169 418
rect 2190 352 2193 478
rect 2206 472 2209 478
rect 2214 462 2217 508
rect 2254 471 2257 558
rect 2250 468 2257 471
rect 2262 462 2265 548
rect 2278 502 2281 538
rect 2278 472 2281 498
rect 2294 472 2297 518
rect 2282 458 2286 461
rect 2214 432 2217 458
rect 2222 452 2225 458
rect 2254 452 2257 458
rect 2198 362 2201 368
rect 2150 288 2158 291
rect 2046 282 2049 288
rect 2118 282 2121 288
rect 2082 278 2089 281
rect 2062 272 2065 278
rect 1974 262 1977 268
rect 1814 252 1817 258
rect 1938 248 1942 251
rect 1926 242 1929 248
rect 1982 242 1985 258
rect 1882 238 1886 241
rect 1994 238 1998 241
rect 1778 218 1782 221
rect 1790 160 1793 179
rect 1846 172 1849 218
rect 1702 152 1705 158
rect 1814 152 1817 158
rect 1742 132 1745 138
rect 1758 122 1761 138
rect 1830 102 1833 138
rect 1750 72 1753 78
rect 1814 72 1817 98
rect 1582 31 1585 50
rect 1446 -18 1449 18
rect 1102 -22 1106 -18
rect 1214 -22 1218 -18
rect 1238 -22 1242 -18
rect 1254 -22 1258 -18
rect 1278 -22 1282 -18
rect 1430 -22 1434 -18
rect 1446 -22 1450 -18
rect 1534 -19 1538 -18
rect 1542 -19 1545 18
rect 1534 -22 1545 -19
rect 1734 -19 1738 -18
rect 1742 -19 1745 18
rect 1734 -22 1745 -19
rect 1862 -18 1865 238
rect 1982 222 1985 238
rect 2006 212 2009 248
rect 2014 212 2017 248
rect 2038 232 2041 268
rect 2078 192 2081 228
rect 1894 132 1897 138
rect 1880 103 1882 107
rect 1886 103 1889 107
rect 1893 103 1896 107
rect 1902 72 1905 188
rect 1918 132 1921 178
rect 1950 160 1953 179
rect 2086 162 2089 278
rect 2102 262 2105 278
rect 2110 272 2113 278
rect 2118 268 2134 271
rect 2118 251 2121 268
rect 2106 248 2121 251
rect 1930 148 1934 151
rect 1982 142 1985 148
rect 2094 142 2097 248
rect 2118 162 2121 168
rect 2102 152 2105 158
rect 2126 142 2129 258
rect 2150 252 2153 278
rect 2166 252 2169 328
rect 2190 261 2193 348
rect 2214 322 2217 348
rect 2214 282 2217 288
rect 2186 258 2193 261
rect 2198 262 2201 278
rect 2206 272 2209 278
rect 2158 152 2161 248
rect 2182 242 2185 248
rect 2190 212 2193 258
rect 2210 248 2214 251
rect 2166 162 2169 208
rect 2198 192 2201 248
rect 2222 242 2225 448
rect 2270 442 2273 458
rect 2230 392 2233 428
rect 2238 382 2241 418
rect 2246 362 2249 368
rect 2230 262 2233 358
rect 2238 342 2241 348
rect 2238 272 2241 278
rect 2246 272 2249 278
rect 2254 262 2257 338
rect 2262 322 2265 348
rect 2270 342 2273 348
rect 2286 342 2289 348
rect 2294 342 2297 468
rect 2302 391 2305 558
rect 2366 542 2369 658
rect 2406 652 2409 658
rect 2384 603 2386 607
rect 2390 603 2393 607
rect 2397 603 2400 607
rect 2430 591 2433 658
rect 2438 602 2441 658
rect 2446 592 2449 668
rect 2470 662 2473 678
rect 2490 668 2494 671
rect 2502 652 2505 658
rect 2474 648 2478 651
rect 2510 642 2513 698
rect 2526 672 2529 768
rect 2566 742 2569 748
rect 2622 742 2625 858
rect 2646 852 2649 858
rect 2654 832 2657 858
rect 2702 842 2705 878
rect 2710 852 2713 1048
rect 2742 1002 2745 1068
rect 2758 1042 2761 1078
rect 2774 1062 2777 1118
rect 2782 1092 2785 1148
rect 2814 1132 2817 1138
rect 2814 1092 2817 1108
rect 2782 1082 2785 1088
rect 2830 1082 2833 1268
rect 2838 1262 2841 1288
rect 2846 1272 2849 1358
rect 2854 1352 2857 1358
rect 2870 1352 2873 1358
rect 2862 1342 2865 1348
rect 2874 1338 2878 1341
rect 2842 1258 2846 1261
rect 2854 1242 2857 1248
rect 2838 1232 2841 1238
rect 2838 1162 2841 1198
rect 2862 1192 2865 1338
rect 2886 1331 2889 1358
rect 2878 1328 2889 1331
rect 2878 1252 2881 1328
rect 2886 1312 2889 1318
rect 2846 1142 2849 1158
rect 2838 1072 2841 1078
rect 2810 1068 2817 1071
rect 2854 1071 2857 1178
rect 2862 1152 2865 1158
rect 2870 1152 2873 1218
rect 2878 1162 2881 1248
rect 2894 1142 2897 1378
rect 2902 1352 2905 1358
rect 2904 1303 2906 1307
rect 2910 1303 2913 1307
rect 2917 1303 2920 1307
rect 2906 1268 2910 1271
rect 2906 1258 2910 1261
rect 2918 1162 2921 1218
rect 2902 1152 2905 1158
rect 2870 1132 2873 1138
rect 2850 1068 2857 1071
rect 2862 1082 2865 1128
rect 2862 1072 2865 1078
rect 2814 1062 2817 1068
rect 2802 1058 2806 1061
rect 2834 1058 2838 1061
rect 2766 1052 2769 1058
rect 2790 1052 2793 1058
rect 2810 1048 2814 1051
rect 2750 1012 2753 1018
rect 2726 962 2729 998
rect 2718 952 2721 958
rect 2774 952 2777 998
rect 2738 948 2742 951
rect 2782 942 2785 968
rect 2726 861 2729 918
rect 2750 872 2753 878
rect 2738 868 2742 871
rect 2726 858 2734 861
rect 2662 792 2665 818
rect 2694 812 2697 818
rect 2702 802 2705 838
rect 2758 822 2761 938
rect 2766 912 2769 918
rect 2790 881 2793 988
rect 2802 958 2814 961
rect 2810 948 2814 951
rect 2798 932 2801 938
rect 2790 878 2801 881
rect 2766 872 2769 878
rect 2798 872 2801 878
rect 2782 862 2785 868
rect 2806 862 2809 938
rect 2830 932 2833 958
rect 2838 952 2841 958
rect 2838 942 2841 948
rect 2846 942 2849 948
rect 2854 941 2857 1068
rect 2862 1042 2865 1048
rect 2886 972 2889 1118
rect 2904 1103 2906 1107
rect 2910 1103 2913 1107
rect 2917 1103 2920 1107
rect 2926 1061 2929 1458
rect 2950 1412 2953 1518
rect 2958 1472 2961 1478
rect 3006 1472 3009 1658
rect 3038 1642 3041 1658
rect 3046 1652 3049 1678
rect 3086 1672 3089 1728
rect 3098 1718 3102 1721
rect 3014 1562 3017 1568
rect 3022 1552 3025 1618
rect 3070 1612 3073 1668
rect 3086 1652 3089 1658
rect 3094 1652 3097 1678
rect 3030 1552 3033 1568
rect 3054 1562 3057 1608
rect 3054 1552 3057 1558
rect 3042 1548 3046 1551
rect 3070 1532 3073 1598
rect 3094 1592 3097 1648
rect 3082 1548 3086 1551
rect 3082 1538 3086 1541
rect 3102 1532 3105 1678
rect 3110 1582 3113 1668
rect 3118 1652 3121 1738
rect 3126 1732 3129 1738
rect 3130 1688 3134 1691
rect 3142 1682 3145 1728
rect 3150 1692 3153 1758
rect 3174 1752 3177 1768
rect 3190 1762 3193 1768
rect 3162 1748 3166 1751
rect 3226 1748 3230 1751
rect 3206 1722 3209 1738
rect 3206 1702 3209 1718
rect 3214 1701 3217 1748
rect 3238 1742 3241 1798
rect 3246 1758 3254 1761
rect 3246 1742 3249 1758
rect 3270 1742 3273 1818
rect 3278 1792 3281 1838
rect 3286 1832 3289 1838
rect 3318 1802 3321 1818
rect 3294 1752 3297 1778
rect 3350 1772 3353 2148
rect 3366 2082 3369 2118
rect 3358 2062 3361 2068
rect 3358 2042 3361 2048
rect 3374 2032 3377 2148
rect 3382 2062 3385 2068
rect 3390 2062 3393 2068
rect 3398 2052 3401 2058
rect 3414 2052 3417 2158
rect 3494 2152 3497 2188
rect 3518 2168 3526 2171
rect 3474 2148 3478 2151
rect 3506 2148 3510 2151
rect 3426 2128 3430 2131
rect 3438 2102 3441 2118
rect 3438 2072 3441 2078
rect 3446 2072 3449 2148
rect 3470 2132 3473 2138
rect 3458 2078 3470 2081
rect 3442 2058 3446 2061
rect 3470 2052 3473 2058
rect 3382 2042 3385 2048
rect 3414 2032 3417 2048
rect 3462 2032 3465 2048
rect 3478 2042 3481 2128
rect 3502 2062 3505 2098
rect 3486 2022 3489 2058
rect 3518 2052 3521 2168
rect 3526 2162 3529 2168
rect 3550 2152 3553 2188
rect 3566 2172 3569 2178
rect 3574 2162 3577 2238
rect 3582 2182 3585 2218
rect 3590 2192 3593 2248
rect 3638 2242 3641 2318
rect 3654 2312 3657 2348
rect 3670 2332 3673 2348
rect 3702 2342 3705 2348
rect 3646 2262 3649 2288
rect 3678 2262 3681 2298
rect 3690 2278 3694 2281
rect 3710 2262 3713 2268
rect 3686 2252 3689 2258
rect 3654 2242 3657 2248
rect 3606 2222 3609 2238
rect 3670 2222 3673 2238
rect 3650 2218 3654 2221
rect 3598 2172 3601 2178
rect 3614 2171 3617 2218
rect 3662 2182 3665 2188
rect 3614 2168 3625 2171
rect 3578 2158 3582 2161
rect 3610 2158 3614 2161
rect 3530 2128 3534 2131
rect 3542 2052 3545 2058
rect 3506 2038 3510 2041
rect 3398 2012 3401 2018
rect 3486 2012 3489 2018
rect 3408 2003 3410 2007
rect 3414 2003 3417 2007
rect 3421 2003 3424 2007
rect 3518 1962 3521 2048
rect 3550 2042 3553 2048
rect 3530 2038 3534 2041
rect 3558 2041 3561 2158
rect 3578 2148 3590 2151
rect 3566 2142 3569 2148
rect 3598 2092 3601 2148
rect 3574 2082 3577 2088
rect 3606 2072 3609 2088
rect 3554 2038 3561 2041
rect 3566 2042 3569 2058
rect 3574 2022 3577 2058
rect 3582 2052 3585 2058
rect 3590 2052 3593 2068
rect 3622 2062 3625 2168
rect 3678 2162 3681 2218
rect 3694 2192 3697 2248
rect 3718 2242 3721 2358
rect 3738 2348 3742 2351
rect 3734 2282 3737 2318
rect 3734 2252 3737 2258
rect 3742 2252 3745 2338
rect 3770 2258 3774 2261
rect 3746 2248 3750 2251
rect 3758 2242 3761 2248
rect 3726 2232 3729 2238
rect 3642 2148 3646 2151
rect 3702 2151 3705 2218
rect 3734 2172 3737 2218
rect 3710 2162 3713 2168
rect 3718 2162 3721 2168
rect 3698 2148 3705 2151
rect 3630 2072 3633 2118
rect 3654 2092 3657 2128
rect 3678 2122 3681 2148
rect 3686 2132 3689 2138
rect 3678 2092 3681 2108
rect 3638 2052 3641 2088
rect 3506 1958 3510 1961
rect 3374 1942 3377 1948
rect 3366 1902 3369 1918
rect 3382 1912 3385 1958
rect 3398 1942 3401 1958
rect 3446 1952 3449 1958
rect 3478 1952 3481 1958
rect 3526 1952 3529 2008
rect 3542 2002 3545 2018
rect 3590 1972 3593 2048
rect 3638 2042 3641 2048
rect 3622 2002 3625 2038
rect 3470 1942 3473 1948
rect 3486 1942 3489 1948
rect 3410 1938 3414 1941
rect 3458 1938 3462 1941
rect 3422 1922 3425 1928
rect 3374 1852 3377 1858
rect 3382 1842 3385 1878
rect 3222 1712 3225 1738
rect 3214 1698 3225 1701
rect 3222 1692 3225 1698
rect 3246 1692 3249 1738
rect 3286 1732 3289 1748
rect 3302 1742 3305 1758
rect 3298 1738 3302 1741
rect 3254 1692 3257 1708
rect 3158 1672 3161 1688
rect 3218 1678 3222 1681
rect 3170 1668 3174 1671
rect 3118 1572 3121 1648
rect 3134 1582 3137 1668
rect 3166 1652 3169 1658
rect 3182 1642 3185 1648
rect 3174 1592 3177 1598
rect 3198 1592 3201 1608
rect 3110 1562 3113 1568
rect 3166 1562 3169 1588
rect 3190 1562 3193 1568
rect 3214 1562 3217 1588
rect 3122 1558 3129 1561
rect 3030 1472 3033 1488
rect 3002 1468 3006 1471
rect 3038 1462 3041 1528
rect 3046 1522 3049 1528
rect 3094 1502 3097 1518
rect 2970 1458 2974 1461
rect 3010 1458 3014 1461
rect 2982 1452 2985 1458
rect 2966 1362 2969 1418
rect 3014 1372 3017 1448
rect 3038 1412 3041 1418
rect 2974 1362 2977 1368
rect 3022 1362 3025 1378
rect 2934 1312 2937 1348
rect 2942 1332 2945 1338
rect 2954 1328 2958 1331
rect 2966 1312 2969 1348
rect 2990 1322 2993 1348
rect 2998 1342 3001 1358
rect 3006 1352 3009 1358
rect 3022 1352 3025 1358
rect 3030 1342 3033 1348
rect 3014 1332 3017 1338
rect 2974 1302 2977 1318
rect 2954 1278 2958 1281
rect 2934 1252 2937 1258
rect 2942 1202 2945 1268
rect 2974 1262 2977 1288
rect 2982 1272 2985 1278
rect 2954 1258 2958 1261
rect 2950 1202 2953 1218
rect 2974 1212 2977 1248
rect 2942 1142 2945 1188
rect 2950 1162 2953 1168
rect 2958 1162 2961 1208
rect 2962 1148 2966 1151
rect 2922 1058 2929 1061
rect 2934 1062 2937 1108
rect 2942 1072 2945 1088
rect 2966 1082 2969 1128
rect 2974 1072 2977 1208
rect 2982 1152 2985 1198
rect 2990 1162 2993 1218
rect 2998 1152 3001 1308
rect 3006 1252 3009 1298
rect 3014 1272 3017 1278
rect 3022 1261 3025 1338
rect 3034 1328 3038 1331
rect 3046 1331 3049 1388
rect 3054 1362 3057 1478
rect 3110 1472 3113 1558
rect 3126 1552 3129 1558
rect 3222 1552 3225 1678
rect 3230 1642 3233 1668
rect 3238 1662 3241 1668
rect 3246 1652 3249 1688
rect 3262 1672 3265 1698
rect 3278 1681 3281 1718
rect 3274 1678 3281 1681
rect 3286 1682 3289 1728
rect 3310 1672 3313 1768
rect 3362 1758 3366 1761
rect 3342 1742 3345 1748
rect 3390 1742 3393 1898
rect 3422 1872 3425 1878
rect 3438 1872 3441 1938
rect 3526 1932 3529 1938
rect 3534 1932 3537 1968
rect 3578 1958 3582 1961
rect 3606 1952 3609 1968
rect 3554 1948 3558 1951
rect 3566 1942 3569 1948
rect 3550 1932 3553 1938
rect 3558 1932 3561 1938
rect 3606 1932 3609 1938
rect 3614 1932 3617 1988
rect 3630 1972 3633 2018
rect 3638 2002 3641 2028
rect 3638 1962 3641 1998
rect 3646 1982 3649 2078
rect 3674 2058 3678 2061
rect 3662 2012 3665 2058
rect 3670 2042 3673 2048
rect 3686 2032 3689 2038
rect 3662 1952 3665 2008
rect 3694 1952 3697 2118
rect 3718 2092 3721 2158
rect 3726 2152 3729 2158
rect 3710 2062 3713 2068
rect 3718 2062 3721 2078
rect 3726 2052 3729 2098
rect 3734 2082 3737 2138
rect 3742 2092 3745 2118
rect 3734 2052 3737 2078
rect 3742 2062 3745 2068
rect 3746 2038 3750 2041
rect 3718 1992 3721 2038
rect 3726 1972 3729 2038
rect 3742 2022 3745 2028
rect 3758 2002 3761 2118
rect 3774 2112 3777 2148
rect 3766 2082 3769 2088
rect 3706 1968 3710 1971
rect 3734 1962 3737 1968
rect 3634 1948 3638 1951
rect 3654 1942 3657 1948
rect 3670 1942 3673 1948
rect 3630 1932 3633 1938
rect 3662 1932 3665 1938
rect 3450 1928 3454 1931
rect 3506 1928 3510 1931
rect 3586 1928 3590 1931
rect 3446 1892 3449 1898
rect 3454 1882 3457 1908
rect 3502 1882 3505 1918
rect 3534 1882 3537 1888
rect 3474 1878 3478 1881
rect 3474 1868 3478 1871
rect 3490 1868 3494 1871
rect 3398 1832 3401 1858
rect 3408 1803 3410 1807
rect 3414 1803 3417 1807
rect 3421 1803 3424 1807
rect 3438 1792 3441 1868
rect 3486 1858 3494 1861
rect 3502 1861 3505 1868
rect 3574 1862 3577 1878
rect 3582 1862 3585 1918
rect 3590 1882 3593 1888
rect 3638 1882 3641 1918
rect 3602 1878 3606 1881
rect 3606 1862 3609 1868
rect 3498 1858 3505 1861
rect 3546 1858 3550 1861
rect 3446 1842 3449 1848
rect 3470 1812 3473 1858
rect 3486 1832 3489 1858
rect 3510 1852 3513 1858
rect 3530 1848 3534 1851
rect 3494 1842 3497 1848
rect 3582 1842 3585 1848
rect 3562 1838 3566 1841
rect 3614 1832 3617 1868
rect 3622 1862 3625 1878
rect 3638 1862 3641 1868
rect 3654 1862 3657 1868
rect 3634 1848 3638 1851
rect 3662 1842 3665 1898
rect 3694 1892 3697 1948
rect 3670 1842 3673 1848
rect 3686 1842 3689 1878
rect 3694 1862 3697 1868
rect 3718 1851 3721 1948
rect 3726 1882 3729 1958
rect 3726 1862 3729 1868
rect 3734 1852 3737 1958
rect 3742 1942 3745 1948
rect 3718 1848 3729 1851
rect 3670 1832 3673 1838
rect 3702 1832 3705 1848
rect 3714 1838 3718 1841
rect 3546 1828 3550 1831
rect 3474 1768 3478 1771
rect 3406 1752 3409 1758
rect 3486 1752 3489 1828
rect 3714 1818 3718 1821
rect 3502 1752 3505 1808
rect 3510 1792 3513 1818
rect 3550 1772 3553 1788
rect 3518 1752 3521 1768
rect 3526 1752 3529 1768
rect 3558 1762 3561 1778
rect 3566 1762 3569 1798
rect 3574 1771 3577 1818
rect 3574 1768 3582 1771
rect 3610 1768 3614 1771
rect 3638 1762 3641 1768
rect 3538 1758 3542 1761
rect 3602 1758 3606 1761
rect 3450 1748 3454 1751
rect 3482 1748 3486 1751
rect 3318 1732 3321 1738
rect 3326 1672 3329 1698
rect 3334 1692 3337 1738
rect 3350 1692 3353 1738
rect 3374 1682 3377 1718
rect 3338 1678 3342 1681
rect 3382 1681 3385 1738
rect 3482 1728 3486 1731
rect 3382 1678 3390 1681
rect 3394 1678 3398 1681
rect 3322 1668 3326 1671
rect 3286 1662 3289 1668
rect 3310 1662 3313 1668
rect 3250 1648 3254 1651
rect 3254 1552 3257 1558
rect 3146 1548 3150 1551
rect 3134 1542 3137 1548
rect 3134 1482 3137 1528
rect 3118 1472 3121 1478
rect 3062 1462 3065 1468
rect 3142 1462 3145 1548
rect 3210 1538 3214 1541
rect 3234 1538 3238 1541
rect 3162 1528 3166 1531
rect 3150 1502 3153 1518
rect 3182 1502 3185 1538
rect 3262 1532 3265 1648
rect 3334 1642 3337 1648
rect 3358 1642 3361 1668
rect 3366 1662 3369 1668
rect 3390 1662 3393 1668
rect 3414 1662 3417 1668
rect 3390 1642 3393 1648
rect 3422 1642 3425 1718
rect 3462 1712 3465 1728
rect 3486 1682 3489 1688
rect 3430 1662 3433 1678
rect 3442 1668 3473 1671
rect 3470 1662 3473 1668
rect 3458 1658 3462 1661
rect 3486 1642 3489 1648
rect 3286 1562 3289 1618
rect 3278 1552 3281 1558
rect 3266 1528 3270 1531
rect 3218 1518 3222 1521
rect 3182 1492 3185 1498
rect 3174 1482 3177 1488
rect 3190 1482 3193 1498
rect 3230 1482 3233 1508
rect 3162 1478 3166 1481
rect 3218 1478 3222 1481
rect 3158 1462 3161 1468
rect 3122 1458 3126 1461
rect 3078 1452 3081 1458
rect 3086 1422 3089 1458
rect 3058 1348 3062 1351
rect 3058 1338 3062 1341
rect 3046 1328 3057 1331
rect 3046 1272 3049 1318
rect 3014 1258 3025 1261
rect 2982 1142 2985 1148
rect 3014 1142 3017 1258
rect 3054 1252 3057 1328
rect 3070 1292 3073 1348
rect 3086 1341 3089 1418
rect 3118 1382 3121 1388
rect 3106 1348 3110 1351
rect 3126 1342 3129 1378
rect 3142 1372 3145 1458
rect 3150 1361 3153 1398
rect 3166 1382 3169 1418
rect 3146 1358 3153 1361
rect 3086 1338 3097 1341
rect 3086 1322 3089 1328
rect 3094 1301 3097 1338
rect 3146 1338 3150 1341
rect 3102 1332 3105 1338
rect 3094 1298 3105 1301
rect 3090 1288 3094 1291
rect 3066 1258 3070 1261
rect 3022 1212 3025 1218
rect 3062 1172 3065 1188
rect 3062 1162 3065 1168
rect 3070 1162 3073 1218
rect 3078 1212 3081 1268
rect 3094 1242 3097 1278
rect 3102 1262 3105 1298
rect 3110 1282 3113 1338
rect 3138 1318 3142 1321
rect 3174 1312 3177 1348
rect 3182 1342 3185 1348
rect 3190 1341 3193 1478
rect 3210 1468 3214 1471
rect 3238 1462 3241 1528
rect 3250 1518 3254 1521
rect 3246 1472 3249 1478
rect 3262 1462 3265 1478
rect 3198 1422 3201 1458
rect 3222 1422 3225 1448
rect 3202 1348 3206 1351
rect 3214 1342 3217 1358
rect 3190 1338 3201 1341
rect 3114 1278 3121 1281
rect 3102 1252 3105 1258
rect 3086 1152 3089 1218
rect 3102 1192 3105 1218
rect 3118 1162 3121 1278
rect 3134 1272 3137 1298
rect 3126 1172 3129 1268
rect 3142 1262 3145 1278
rect 3166 1272 3169 1298
rect 3182 1261 3185 1338
rect 3198 1332 3201 1338
rect 3190 1302 3193 1318
rect 3222 1312 3225 1418
rect 3230 1342 3233 1348
rect 3238 1342 3241 1408
rect 3254 1372 3257 1458
rect 3254 1362 3257 1368
rect 3258 1348 3262 1351
rect 3230 1322 3233 1328
rect 3214 1282 3217 1288
rect 3230 1282 3233 1298
rect 3238 1282 3241 1338
rect 3270 1272 3273 1518
rect 3278 1332 3281 1548
rect 3286 1542 3289 1548
rect 3294 1542 3297 1588
rect 3310 1572 3313 1618
rect 3408 1603 3410 1607
rect 3414 1603 3417 1607
rect 3421 1603 3424 1607
rect 3318 1552 3321 1558
rect 3358 1552 3361 1558
rect 3310 1532 3313 1538
rect 3318 1532 3321 1548
rect 3350 1542 3353 1548
rect 3366 1542 3369 1578
rect 3390 1552 3393 1568
rect 3398 1552 3401 1578
rect 3374 1542 3377 1548
rect 3422 1542 3425 1568
rect 3454 1552 3457 1588
rect 3402 1538 3406 1541
rect 3306 1518 3310 1521
rect 3310 1508 3318 1511
rect 3286 1472 3289 1508
rect 3294 1482 3297 1508
rect 3298 1468 3302 1471
rect 3294 1422 3297 1458
rect 3298 1358 3302 1361
rect 3278 1272 3281 1318
rect 3294 1292 3297 1338
rect 3286 1272 3289 1288
rect 3302 1282 3305 1328
rect 3310 1292 3313 1508
rect 3326 1502 3329 1528
rect 3342 1522 3345 1538
rect 3334 1511 3337 1518
rect 3334 1508 3342 1511
rect 3366 1462 3369 1468
rect 3358 1452 3361 1458
rect 3326 1392 3329 1438
rect 3318 1342 3321 1348
rect 3334 1342 3337 1428
rect 3342 1372 3345 1418
rect 3342 1342 3345 1348
rect 3350 1342 3353 1348
rect 3370 1338 3374 1341
rect 3350 1292 3353 1338
rect 3362 1328 3366 1331
rect 3358 1312 3361 1318
rect 3382 1302 3385 1538
rect 3398 1482 3401 1488
rect 3414 1472 3417 1538
rect 3430 1522 3433 1548
rect 3462 1542 3465 1638
rect 3494 1622 3497 1678
rect 3502 1662 3505 1748
rect 3514 1658 3518 1661
rect 3526 1652 3529 1658
rect 3534 1651 3537 1758
rect 3566 1752 3569 1758
rect 3590 1752 3593 1758
rect 3630 1752 3633 1758
rect 3646 1752 3649 1818
rect 3554 1748 3558 1751
rect 3542 1692 3545 1748
rect 3590 1732 3593 1738
rect 3574 1682 3577 1708
rect 3546 1678 3550 1681
rect 3566 1672 3569 1678
rect 3598 1672 3601 1678
rect 3614 1672 3617 1748
rect 3630 1682 3633 1698
rect 3590 1662 3593 1668
rect 3570 1658 3574 1661
rect 3534 1648 3542 1651
rect 3598 1651 3601 1658
rect 3590 1648 3601 1651
rect 3534 1642 3537 1648
rect 3590 1642 3593 1648
rect 3470 1542 3473 1548
rect 3390 1362 3393 1468
rect 3422 1462 3425 1518
rect 3446 1432 3449 1468
rect 3454 1462 3457 1478
rect 3402 1418 3406 1421
rect 3408 1403 3410 1407
rect 3414 1403 3417 1407
rect 3421 1403 3424 1407
rect 3398 1352 3401 1388
rect 3454 1362 3457 1418
rect 3470 1392 3473 1518
rect 3478 1482 3481 1578
rect 3494 1562 3497 1598
rect 3502 1582 3505 1628
rect 3622 1602 3625 1648
rect 3638 1592 3641 1698
rect 3654 1682 3657 1778
rect 3662 1772 3665 1778
rect 3674 1768 3678 1771
rect 3694 1771 3697 1818
rect 3694 1768 3705 1771
rect 3678 1742 3681 1758
rect 3694 1752 3697 1758
rect 3686 1732 3689 1748
rect 3670 1702 3673 1718
rect 3646 1672 3649 1678
rect 3678 1672 3681 1678
rect 3694 1672 3697 1738
rect 3702 1672 3705 1768
rect 3670 1662 3673 1668
rect 3658 1658 3662 1661
rect 3682 1658 3686 1661
rect 3646 1632 3649 1658
rect 3694 1652 3697 1658
rect 3670 1592 3673 1628
rect 3702 1602 3705 1648
rect 3710 1622 3713 1768
rect 3718 1752 3721 1758
rect 3726 1731 3729 1848
rect 3734 1752 3737 1848
rect 3742 1842 3745 1918
rect 3754 1858 3758 1861
rect 3766 1852 3769 1878
rect 3754 1838 3758 1841
rect 3742 1802 3745 1818
rect 3750 1768 3758 1771
rect 3742 1762 3745 1768
rect 3750 1751 3753 1768
rect 3766 1762 3769 1848
rect 3774 1792 3777 2018
rect 3770 1758 3774 1761
rect 3742 1748 3753 1751
rect 3762 1748 3766 1751
rect 3734 1742 3737 1748
rect 3726 1728 3737 1731
rect 3718 1662 3721 1718
rect 3726 1662 3729 1688
rect 3734 1681 3737 1728
rect 3742 1692 3745 1748
rect 3750 1712 3753 1718
rect 3734 1678 3745 1681
rect 3718 1642 3721 1648
rect 3726 1632 3729 1648
rect 3734 1642 3737 1648
rect 3742 1632 3745 1678
rect 3754 1658 3758 1661
rect 3766 1652 3769 1718
rect 3750 1648 3758 1651
rect 3750 1642 3753 1648
rect 3538 1588 3542 1591
rect 3490 1548 3494 1551
rect 3486 1532 3489 1538
rect 3494 1502 3497 1518
rect 3450 1348 3454 1351
rect 3406 1342 3409 1348
rect 3406 1322 3409 1338
rect 3418 1328 3422 1331
rect 3358 1282 3361 1288
rect 3342 1272 3345 1278
rect 3242 1268 3246 1271
rect 3322 1268 3326 1271
rect 3182 1258 3190 1261
rect 3242 1258 3246 1261
rect 3042 1148 3046 1151
rect 3058 1138 3062 1141
rect 2986 1128 2990 1131
rect 2998 1121 3001 1138
rect 3006 1132 3009 1138
rect 3030 1132 3033 1138
rect 3038 1132 3041 1138
rect 3066 1128 3070 1131
rect 2998 1118 3006 1121
rect 3026 1118 3030 1121
rect 3022 1092 3025 1108
rect 3042 1078 3054 1081
rect 3074 1078 3078 1081
rect 2974 1062 2977 1068
rect 2954 1058 2958 1061
rect 3058 1058 3062 1061
rect 2998 1052 3001 1058
rect 2918 1022 2921 1048
rect 2934 1032 2937 1038
rect 3014 1022 3017 1048
rect 2934 992 2937 1018
rect 2950 1002 2953 1018
rect 2990 1002 2993 1018
rect 2958 962 2961 968
rect 3014 962 3017 968
rect 2906 958 2910 961
rect 2946 958 2950 961
rect 2882 948 2886 951
rect 2922 948 2926 951
rect 2978 948 2982 951
rect 3002 948 3006 951
rect 2854 938 2862 941
rect 2850 928 2854 931
rect 2814 872 2817 918
rect 2830 902 2833 918
rect 2870 912 2873 948
rect 2878 901 2881 938
rect 2926 932 2929 938
rect 2904 903 2906 907
rect 2910 903 2913 907
rect 2917 903 2920 907
rect 2870 898 2881 901
rect 2846 872 2849 878
rect 2870 872 2873 898
rect 2882 878 2886 881
rect 2922 878 2926 881
rect 2934 872 2937 948
rect 2990 942 2993 948
rect 2962 918 2969 921
rect 2958 882 2961 908
rect 2958 872 2961 878
rect 2966 872 2969 918
rect 2982 882 2985 938
rect 2990 872 2993 918
rect 2770 858 2774 861
rect 2818 858 2822 861
rect 2838 852 2841 868
rect 2766 842 2769 848
rect 2802 838 2806 841
rect 2702 752 2705 768
rect 2734 752 2737 818
rect 2762 748 2766 751
rect 2694 742 2697 748
rect 2726 742 2729 748
rect 2750 742 2753 748
rect 2738 738 2742 741
rect 2774 732 2777 798
rect 2798 752 2801 768
rect 2822 752 2825 818
rect 2846 792 2849 868
rect 2854 842 2857 858
rect 2894 842 2897 868
rect 2902 862 2905 868
rect 2934 842 2937 848
rect 2854 772 2857 818
rect 2862 772 2865 778
rect 2674 728 2678 731
rect 2722 728 2726 731
rect 2538 688 2542 691
rect 2430 588 2441 591
rect 2414 562 2417 588
rect 2438 552 2441 588
rect 2450 558 2454 561
rect 2350 532 2353 538
rect 2390 492 2393 498
rect 2314 478 2318 481
rect 2310 462 2313 468
rect 2326 462 2329 488
rect 2334 472 2337 478
rect 2366 462 2369 478
rect 2374 462 2377 468
rect 2342 452 2345 458
rect 2310 422 2313 428
rect 2350 401 2353 448
rect 2346 398 2353 401
rect 2302 388 2313 391
rect 2310 362 2313 388
rect 2342 362 2345 398
rect 2314 358 2318 361
rect 2338 348 2342 351
rect 2302 342 2305 348
rect 2338 338 2342 341
rect 2358 341 2361 458
rect 2382 442 2385 468
rect 2366 382 2369 418
rect 2374 382 2377 408
rect 2384 403 2386 407
rect 2390 403 2393 407
rect 2397 403 2400 407
rect 2374 362 2377 378
rect 2398 352 2401 358
rect 2366 342 2369 348
rect 2358 338 2366 341
rect 2282 328 2310 331
rect 2286 272 2289 308
rect 2342 292 2345 328
rect 2298 288 2302 291
rect 2270 242 2273 248
rect 2182 162 2185 188
rect 2198 158 2206 161
rect 2166 152 2169 158
rect 2190 152 2193 158
rect 2138 148 2142 151
rect 2150 142 2153 148
rect 2158 142 2161 148
rect 2182 142 2185 148
rect 1918 82 1921 128
rect 1998 102 2001 128
rect 2126 122 2129 128
rect 2006 82 2009 108
rect 2094 82 2097 88
rect 2078 72 2081 78
rect 2179 68 2182 71
rect 2038 62 2041 68
rect 2134 62 2137 68
rect 1962 58 1966 61
rect 2190 52 2193 148
rect 2198 92 2201 158
rect 2230 152 2233 208
rect 2242 158 2246 161
rect 2254 151 2257 218
rect 2254 148 2262 151
rect 2206 142 2209 148
rect 2270 142 2273 198
rect 2278 172 2281 258
rect 2278 152 2281 168
rect 2234 138 2238 141
rect 2250 138 2254 141
rect 2206 112 2209 138
rect 2214 92 2217 118
rect 2210 68 2214 71
rect 2230 62 2233 108
rect 2278 72 2281 118
rect 2294 112 2297 148
rect 2302 102 2305 268
rect 2310 222 2313 258
rect 2350 212 2353 338
rect 2310 160 2313 179
rect 2358 162 2361 278
rect 2382 262 2385 328
rect 2390 302 2393 348
rect 2406 332 2409 548
rect 2454 502 2457 558
rect 2454 482 2457 488
rect 2414 472 2417 478
rect 2462 472 2465 548
rect 2470 492 2473 548
rect 2486 541 2489 638
rect 2482 538 2489 541
rect 2478 482 2481 488
rect 2486 482 2489 518
rect 2494 472 2497 608
rect 2582 602 2585 728
rect 2662 702 2665 718
rect 2686 682 2689 718
rect 2710 682 2713 728
rect 2726 682 2729 698
rect 2622 612 2625 678
rect 2638 672 2641 678
rect 2734 672 2737 688
rect 2750 672 2753 698
rect 2798 692 2801 738
rect 2810 728 2814 731
rect 2814 712 2817 718
rect 2822 682 2825 748
rect 2830 742 2833 748
rect 2838 742 2841 768
rect 2886 762 2889 798
rect 2910 762 2913 768
rect 2886 752 2889 758
rect 2922 748 2926 751
rect 2878 742 2881 748
rect 2934 742 2937 788
rect 2854 732 2857 738
rect 2862 732 2865 738
rect 2942 732 2945 868
rect 2986 858 2990 861
rect 2950 812 2953 858
rect 2966 842 2969 848
rect 2974 782 2977 858
rect 2998 852 3001 938
rect 3022 922 3025 1028
rect 3030 961 3033 1028
rect 3050 1018 3054 1021
rect 3050 978 3054 981
rect 3038 972 3041 978
rect 3030 958 3041 961
rect 3030 932 3033 948
rect 3038 882 3041 958
rect 3070 952 3073 1048
rect 3078 982 3081 1058
rect 3078 962 3081 968
rect 3086 952 3089 1128
rect 3094 1092 3097 1138
rect 3102 1112 3105 1148
rect 3118 1112 3121 1148
rect 3126 1142 3129 1168
rect 3134 1152 3137 1158
rect 3126 1092 3129 1118
rect 3118 1072 3121 1088
rect 3142 1082 3145 1248
rect 3158 1162 3161 1248
rect 3154 1158 3158 1161
rect 3166 1151 3169 1198
rect 3162 1148 3169 1151
rect 3158 1142 3161 1148
rect 3166 1132 3169 1138
rect 3142 1072 3145 1078
rect 3150 1062 3153 1068
rect 3106 1058 3110 1061
rect 3094 1052 3097 1058
rect 3142 1052 3145 1058
rect 3106 1048 3110 1051
rect 3098 1038 3102 1041
rect 3134 952 3137 1038
rect 3150 962 3153 968
rect 3142 952 3145 958
rect 3058 948 3062 951
rect 3130 948 3134 951
rect 3118 942 3121 948
rect 3030 872 3033 878
rect 3046 872 3049 888
rect 3014 862 3017 868
rect 2938 728 2942 731
rect 2846 711 2849 718
rect 2846 708 2857 711
rect 2838 692 2841 708
rect 2762 678 2766 681
rect 2778 668 2782 671
rect 2710 662 2713 668
rect 2670 631 2673 650
rect 2522 588 2526 591
rect 2670 562 2673 588
rect 2678 552 2681 658
rect 2690 558 2694 561
rect 2714 558 2718 561
rect 2726 552 2729 598
rect 2506 548 2510 551
rect 2706 548 2710 551
rect 2622 542 2625 548
rect 2522 538 2526 541
rect 2606 522 2609 528
rect 2558 492 2561 518
rect 2622 511 2625 518
rect 2614 508 2625 511
rect 2614 492 2617 508
rect 2654 482 2657 548
rect 2718 542 2721 548
rect 2734 542 2737 668
rect 2790 662 2793 668
rect 2746 658 2750 661
rect 2782 642 2785 658
rect 2830 642 2833 668
rect 2838 651 2841 678
rect 2846 672 2849 698
rect 2854 692 2857 708
rect 2894 702 2897 718
rect 2904 703 2906 707
rect 2910 703 2913 707
rect 2917 703 2920 707
rect 2874 688 2878 691
rect 2906 688 2910 691
rect 2882 668 2886 671
rect 2850 658 2854 661
rect 2838 648 2846 651
rect 2886 642 2889 658
rect 2894 652 2897 688
rect 2950 682 2953 778
rect 2958 752 2961 768
rect 2974 762 2977 768
rect 2978 748 2985 751
rect 2962 738 2966 741
rect 2982 732 2985 748
rect 2998 742 3001 848
rect 3006 792 3009 818
rect 3022 772 3025 868
rect 3054 842 3057 938
rect 3070 852 3073 938
rect 3086 862 3089 918
rect 3094 882 3097 938
rect 3134 932 3137 938
rect 3114 928 3118 931
rect 3102 902 3105 918
rect 3126 872 3129 888
rect 3142 872 3145 948
rect 3098 868 3102 871
rect 3114 858 3118 861
rect 3030 752 3033 768
rect 3018 748 3022 751
rect 3014 732 3017 738
rect 2962 728 2966 731
rect 2982 692 2985 728
rect 2930 678 2934 681
rect 2910 642 2913 668
rect 2950 662 2953 678
rect 2974 662 2977 668
rect 2990 661 2993 698
rect 2998 682 3001 728
rect 3022 672 3025 738
rect 3030 681 3033 748
rect 3046 732 3049 808
rect 3062 742 3065 818
rect 3054 732 3057 738
rect 3038 712 3041 718
rect 3030 678 3038 681
rect 3006 662 3009 668
rect 3062 662 3065 718
rect 3070 692 3073 838
rect 3086 832 3089 838
rect 3102 822 3105 848
rect 3118 842 3121 848
rect 3094 772 3097 778
rect 3078 762 3081 768
rect 3102 742 3105 818
rect 3134 792 3137 868
rect 3142 832 3145 858
rect 3142 781 3145 818
rect 3150 812 3153 918
rect 3158 902 3161 1128
rect 3166 1092 3169 1118
rect 3174 1002 3177 1218
rect 3182 1202 3185 1258
rect 3190 1222 3193 1248
rect 3202 1238 3206 1241
rect 3222 1202 3225 1218
rect 3218 1188 3222 1191
rect 3270 1182 3273 1268
rect 3278 1172 3281 1258
rect 3306 1248 3310 1251
rect 3286 1192 3289 1248
rect 3334 1232 3337 1258
rect 3182 1112 3185 1168
rect 3342 1162 3345 1268
rect 3374 1262 3377 1268
rect 3390 1252 3393 1318
rect 3414 1312 3417 1318
rect 3398 1272 3401 1308
rect 3422 1282 3425 1328
rect 3454 1272 3457 1308
rect 3462 1292 3465 1368
rect 3478 1332 3481 1478
rect 3494 1472 3497 1478
rect 3502 1462 3505 1578
rect 3514 1548 3518 1551
rect 3526 1542 3529 1568
rect 3534 1531 3537 1558
rect 3542 1552 3545 1568
rect 3554 1558 3558 1561
rect 3574 1551 3577 1568
rect 3622 1562 3625 1568
rect 3586 1558 3590 1561
rect 3574 1548 3582 1551
rect 3610 1548 3614 1551
rect 3638 1542 3641 1548
rect 3610 1538 3614 1541
rect 3530 1528 3542 1531
rect 3538 1478 3542 1481
rect 3550 1471 3553 1518
rect 3574 1512 3577 1518
rect 3542 1468 3553 1471
rect 3558 1472 3561 1478
rect 3530 1458 3534 1461
rect 3502 1352 3505 1448
rect 3542 1392 3545 1468
rect 3582 1462 3585 1498
rect 3590 1492 3593 1518
rect 3614 1492 3617 1528
rect 3622 1522 3625 1528
rect 3638 1522 3641 1528
rect 3590 1462 3593 1468
rect 3550 1452 3553 1458
rect 3558 1452 3561 1458
rect 3614 1452 3617 1478
rect 3558 1381 3561 1448
rect 3622 1442 3625 1478
rect 3630 1461 3633 1498
rect 3646 1482 3649 1578
rect 3694 1568 3702 1571
rect 3654 1532 3657 1558
rect 3682 1548 3686 1551
rect 3670 1502 3673 1518
rect 3694 1492 3697 1568
rect 3734 1562 3737 1568
rect 3722 1558 3726 1561
rect 3710 1532 3713 1548
rect 3702 1492 3705 1518
rect 3658 1478 3662 1481
rect 3642 1468 3646 1471
rect 3666 1468 3670 1471
rect 3678 1462 3681 1478
rect 3630 1458 3638 1461
rect 3662 1452 3665 1458
rect 3550 1378 3561 1381
rect 3550 1362 3553 1378
rect 3558 1362 3561 1368
rect 3526 1342 3529 1348
rect 3542 1342 3545 1348
rect 3550 1341 3553 1358
rect 3566 1352 3569 1378
rect 3646 1362 3649 1428
rect 3602 1348 3606 1351
rect 3626 1348 3630 1351
rect 3650 1348 3654 1351
rect 3566 1342 3569 1348
rect 3574 1342 3577 1348
rect 3550 1338 3561 1341
rect 3618 1338 3622 1341
rect 3650 1338 3654 1341
rect 3478 1292 3481 1328
rect 3510 1322 3513 1328
rect 3522 1318 3526 1321
rect 3418 1268 3422 1271
rect 3474 1268 3478 1271
rect 3406 1252 3409 1268
rect 3422 1222 3425 1268
rect 3446 1252 3449 1258
rect 3366 1182 3369 1188
rect 3374 1172 3377 1218
rect 3408 1203 3410 1207
rect 3414 1203 3417 1207
rect 3421 1203 3424 1207
rect 3478 1181 3481 1258
rect 3486 1252 3489 1318
rect 3534 1312 3537 1338
rect 3550 1292 3553 1308
rect 3542 1272 3545 1288
rect 3558 1282 3561 1338
rect 3598 1332 3601 1338
rect 3586 1328 3590 1331
rect 3618 1328 3622 1331
rect 3582 1312 3585 1318
rect 3646 1292 3649 1298
rect 3578 1288 3582 1291
rect 3602 1288 3606 1291
rect 3494 1262 3497 1268
rect 3502 1242 3505 1268
rect 3486 1192 3489 1208
rect 3510 1192 3513 1268
rect 3530 1248 3534 1251
rect 3550 1182 3553 1188
rect 3478 1178 3489 1181
rect 3322 1158 3326 1161
rect 3474 1158 3478 1161
rect 3206 1152 3209 1158
rect 3190 1132 3193 1138
rect 3182 1062 3185 1108
rect 3182 942 3185 968
rect 3190 942 3193 1078
rect 3222 1072 3225 1148
rect 3230 1132 3233 1148
rect 3238 1142 3241 1148
rect 3246 1132 3249 1148
rect 3254 1142 3257 1158
rect 3370 1148 3374 1151
rect 3450 1148 3454 1151
rect 3330 1138 3334 1141
rect 3274 1128 3278 1131
rect 3230 1102 3233 1128
rect 3286 1121 3289 1138
rect 3278 1118 3289 1121
rect 3302 1122 3305 1138
rect 3246 1092 3249 1118
rect 3278 1092 3281 1118
rect 3334 1082 3337 1088
rect 3250 1078 3254 1081
rect 3342 1072 3345 1148
rect 3350 1142 3353 1148
rect 3386 1128 3390 1131
rect 3358 1072 3361 1078
rect 3222 1062 3225 1068
rect 3238 1062 3241 1068
rect 3210 1058 3214 1061
rect 3230 1052 3233 1058
rect 3262 1032 3265 1068
rect 3286 1062 3289 1068
rect 3314 1058 3318 1061
rect 3282 1048 3286 1051
rect 3294 1032 3297 1058
rect 3342 1032 3345 1068
rect 3406 1062 3409 1148
rect 3462 1142 3465 1148
rect 3478 1142 3481 1148
rect 3446 1132 3449 1138
rect 3454 1132 3457 1138
rect 3486 1132 3489 1178
rect 3494 1172 3497 1178
rect 3534 1161 3537 1168
rect 3534 1158 3545 1161
rect 3418 1128 3422 1131
rect 3430 1122 3433 1128
rect 3438 1092 3441 1108
rect 3470 1092 3473 1128
rect 3494 1122 3497 1148
rect 3502 1111 3505 1158
rect 3542 1152 3545 1158
rect 3530 1148 3534 1151
rect 3514 1128 3518 1131
rect 3494 1108 3505 1111
rect 3430 1072 3433 1078
rect 3462 1072 3465 1088
rect 3474 1078 3478 1081
rect 3378 1058 3382 1061
rect 3442 1058 3446 1061
rect 3350 1042 3353 1048
rect 3202 1018 3206 1021
rect 3202 958 3206 961
rect 3170 938 3174 941
rect 3170 928 3174 931
rect 3166 872 3169 888
rect 3170 858 3174 861
rect 3182 851 3185 938
rect 3214 932 3217 1028
rect 3310 992 3313 1018
rect 3230 952 3233 958
rect 3262 952 3265 958
rect 3290 948 3294 951
rect 3206 882 3209 918
rect 3202 868 3206 871
rect 3214 862 3217 928
rect 3230 862 3233 898
rect 3238 862 3241 938
rect 3246 932 3249 948
rect 3298 938 3302 941
rect 3266 928 3270 931
rect 3262 881 3265 918
rect 3278 882 3281 938
rect 3286 932 3289 938
rect 3294 912 3297 928
rect 3302 882 3305 888
rect 3262 878 3270 881
rect 3266 868 3270 871
rect 3246 862 3249 868
rect 3254 852 3257 868
rect 3286 858 3294 861
rect 3182 848 3190 851
rect 3158 842 3161 848
rect 3174 842 3177 848
rect 3182 822 3185 848
rect 3142 778 3153 781
rect 3110 752 3113 758
rect 3134 742 3137 758
rect 3142 752 3145 768
rect 3086 732 3089 738
rect 3118 732 3121 738
rect 3134 722 3137 728
rect 3106 688 3110 691
rect 3078 672 3081 688
rect 3098 668 3102 671
rect 2982 658 2993 661
rect 3034 658 3046 661
rect 2974 642 2977 648
rect 2742 602 2745 618
rect 2742 552 2745 598
rect 2758 592 2761 638
rect 2766 562 2769 568
rect 2798 562 2801 568
rect 2822 562 2825 638
rect 2942 612 2945 618
rect 2866 558 2870 561
rect 2766 542 2769 558
rect 2878 552 2881 598
rect 2886 552 2889 568
rect 2942 552 2945 558
rect 2778 548 2782 551
rect 2866 548 2870 551
rect 2914 548 2918 551
rect 2886 542 2889 548
rect 2794 538 2798 541
rect 2810 538 2814 541
rect 2958 541 2961 568
rect 2966 552 2969 558
rect 2974 542 2977 548
rect 2958 538 2966 541
rect 2498 468 2502 471
rect 2594 468 2598 471
rect 2446 462 2449 468
rect 2434 458 2438 461
rect 2458 458 2462 461
rect 2414 392 2417 458
rect 2438 432 2441 448
rect 2422 392 2425 398
rect 2446 392 2449 458
rect 2486 441 2489 468
rect 2498 458 2502 461
rect 2574 442 2577 468
rect 2590 442 2593 458
rect 2486 438 2494 441
rect 2462 362 2465 388
rect 2502 361 2505 428
rect 2514 368 2518 371
rect 2502 358 2513 361
rect 2414 342 2417 358
rect 2438 352 2441 358
rect 2426 338 2430 341
rect 2454 331 2457 358
rect 2462 352 2465 358
rect 2494 352 2497 358
rect 2470 342 2473 348
rect 2502 342 2505 348
rect 2510 342 2513 358
rect 2454 328 2470 331
rect 2422 282 2425 328
rect 2438 272 2441 288
rect 2478 252 2481 318
rect 2510 292 2513 338
rect 2526 272 2529 418
rect 2534 262 2537 438
rect 2614 432 2617 468
rect 2626 458 2630 461
rect 2630 442 2633 448
rect 2558 402 2561 418
rect 2582 412 2585 418
rect 2582 392 2585 408
rect 2590 332 2593 398
rect 2606 342 2609 398
rect 2638 352 2641 478
rect 2662 472 2665 478
rect 2650 468 2654 471
rect 2646 442 2649 458
rect 2654 431 2657 458
rect 2694 452 2697 538
rect 2718 472 2721 478
rect 2742 472 2745 518
rect 2750 472 2753 528
rect 2774 472 2777 538
rect 2822 532 2825 538
rect 2834 528 2838 531
rect 2818 518 2822 521
rect 2710 462 2713 468
rect 2746 458 2750 461
rect 2758 452 2761 458
rect 2714 448 2726 451
rect 2686 442 2689 448
rect 2650 428 2657 431
rect 2654 362 2657 388
rect 2670 352 2673 418
rect 2694 372 2697 448
rect 2742 402 2745 418
rect 2742 362 2745 388
rect 2762 368 2766 371
rect 2706 358 2710 361
rect 2698 348 2702 351
rect 2722 348 2726 351
rect 2542 272 2545 308
rect 2550 292 2553 298
rect 2558 272 2561 308
rect 2470 231 2473 250
rect 2384 203 2386 207
rect 2390 203 2393 207
rect 2397 203 2400 207
rect 2434 188 2438 191
rect 2474 188 2478 191
rect 2486 162 2489 258
rect 2506 248 2510 251
rect 2534 232 2537 258
rect 2558 212 2561 268
rect 2566 262 2569 298
rect 2582 272 2585 308
rect 2590 282 2593 328
rect 2622 292 2625 298
rect 2594 268 2598 271
rect 2574 262 2577 268
rect 2614 262 2617 278
rect 2654 262 2657 348
rect 2734 342 2737 358
rect 2766 352 2769 358
rect 2774 352 2777 468
rect 2782 392 2785 468
rect 2790 452 2793 498
rect 2814 472 2817 498
rect 2830 492 2833 498
rect 2846 492 2849 538
rect 2918 532 2921 538
rect 2866 528 2870 531
rect 2822 472 2825 488
rect 2870 472 2873 478
rect 2842 468 2846 471
rect 2802 448 2806 451
rect 2814 422 2817 458
rect 2822 442 2825 468
rect 2874 458 2878 461
rect 2838 452 2841 458
rect 2854 451 2857 458
rect 2850 448 2857 451
rect 2866 448 2870 451
rect 2754 348 2758 351
rect 2698 338 2702 341
rect 2714 338 2718 341
rect 2762 338 2766 341
rect 2678 302 2681 328
rect 2686 302 2689 318
rect 2702 272 2705 298
rect 2590 252 2593 258
rect 2342 142 2345 148
rect 2358 132 2361 158
rect 2398 152 2401 158
rect 2518 152 2521 158
rect 2574 142 2577 198
rect 2558 132 2561 138
rect 2606 102 2609 258
rect 2630 242 2633 258
rect 2622 162 2625 188
rect 2630 152 2633 188
rect 2646 132 2649 228
rect 2654 192 2657 258
rect 2662 152 2665 238
rect 2670 231 2673 250
rect 2718 182 2721 278
rect 2774 222 2777 338
rect 2742 182 2745 188
rect 2706 158 2710 161
rect 2722 148 2726 151
rect 2690 138 2694 141
rect 2730 138 2734 141
rect 2646 112 2649 128
rect 2678 122 2681 128
rect 2294 82 2297 98
rect 2374 92 2377 98
rect 2586 88 2590 91
rect 2294 72 2297 78
rect 2494 72 2497 78
rect 2670 72 2673 78
rect 2758 72 2761 78
rect 2510 62 2513 68
rect 2630 62 2633 68
rect 2686 62 2689 68
rect 2782 62 2785 388
rect 2798 352 2801 368
rect 2818 358 2822 361
rect 2790 342 2793 348
rect 2830 341 2833 368
rect 2862 362 2865 448
rect 2854 352 2857 358
rect 2878 352 2881 458
rect 2894 452 2897 518
rect 2904 503 2906 507
rect 2910 503 2913 507
rect 2917 503 2920 507
rect 2926 471 2929 518
rect 2918 468 2929 471
rect 2942 472 2945 478
rect 2974 472 2977 538
rect 2982 472 2985 658
rect 2990 642 2993 648
rect 2990 562 2993 638
rect 2998 542 3001 658
rect 3014 642 3017 658
rect 3062 642 3065 648
rect 3054 562 3057 618
rect 3018 558 3022 561
rect 3030 552 3033 558
rect 3010 548 3014 551
rect 3054 542 3057 558
rect 3070 542 3073 548
rect 3002 538 3006 541
rect 3022 512 3025 518
rect 3038 502 3041 538
rect 3058 528 3062 531
rect 3078 522 3081 658
rect 3110 632 3113 668
rect 3118 662 3121 668
rect 3126 662 3129 718
rect 3110 582 3113 628
rect 3090 558 3094 561
rect 3118 552 3121 568
rect 3126 552 3129 658
rect 3142 622 3145 638
rect 3142 562 3145 618
rect 3086 532 3089 538
rect 3046 482 3049 518
rect 2894 442 2897 448
rect 2894 392 2897 398
rect 2910 342 2913 468
rect 2918 372 2921 468
rect 2930 458 2934 461
rect 2942 458 2950 461
rect 2970 458 2974 461
rect 3026 458 3030 461
rect 2942 452 2945 458
rect 2950 452 2953 458
rect 2990 452 2993 458
rect 2934 362 2937 418
rect 2942 362 2945 448
rect 2966 442 2969 448
rect 3014 432 3017 448
rect 2990 401 2993 418
rect 2982 398 2993 401
rect 2966 362 2969 388
rect 2974 372 2977 388
rect 2982 382 2985 398
rect 3038 392 3041 468
rect 3050 448 3054 451
rect 2974 352 2977 368
rect 2922 348 2926 351
rect 3014 342 3017 358
rect 2826 338 2833 341
rect 2822 292 2825 328
rect 2878 322 2881 338
rect 2886 332 2889 338
rect 2846 272 2849 318
rect 2854 272 2857 318
rect 2904 303 2906 307
rect 2910 303 2913 307
rect 2917 303 2920 307
rect 2862 272 2865 278
rect 2794 258 2799 261
rect 2842 258 2846 261
rect 2830 222 2833 248
rect 2846 242 2849 248
rect 2830 152 2833 168
rect 2838 142 2841 238
rect 2854 192 2857 268
rect 2870 262 2873 298
rect 2934 291 2937 338
rect 2926 288 2937 291
rect 2898 248 2902 251
rect 2886 242 2889 248
rect 2874 218 2878 221
rect 2846 142 2849 148
rect 2798 132 2801 138
rect 2822 72 2825 128
rect 2838 101 2841 138
rect 2830 98 2841 101
rect 2830 62 2833 98
rect 2846 91 2849 118
rect 2842 88 2849 91
rect 2854 92 2857 98
rect 2854 82 2857 88
rect 2870 82 2873 208
rect 2882 148 2886 151
rect 2886 72 2889 78
rect 2894 72 2897 218
rect 2910 202 2913 268
rect 2926 262 2929 288
rect 2938 278 2942 281
rect 2950 271 2953 308
rect 2946 268 2953 271
rect 2958 272 2961 328
rect 2982 272 2985 278
rect 2934 152 2937 258
rect 2942 242 2945 248
rect 2974 232 2977 268
rect 2990 252 2993 298
rect 3014 272 3017 278
rect 3022 262 3025 268
rect 3010 258 3014 261
rect 3018 248 3022 251
rect 2958 162 2961 168
rect 2946 158 2950 161
rect 2974 152 2977 178
rect 2962 148 2966 151
rect 2926 142 2929 148
rect 2982 142 2985 228
rect 3006 192 3009 218
rect 3030 202 3033 328
rect 3038 262 3041 288
rect 3070 272 3073 498
rect 3078 392 3081 518
rect 3094 462 3097 538
rect 3142 532 3145 538
rect 3134 482 3137 488
rect 3150 472 3153 778
rect 3186 768 3190 771
rect 3170 758 3174 761
rect 3190 742 3193 748
rect 3206 742 3209 848
rect 3214 842 3217 848
rect 3230 792 3233 818
rect 3230 742 3233 768
rect 3238 752 3241 838
rect 3258 758 3262 761
rect 3286 752 3289 858
rect 3310 841 3313 948
rect 3318 932 3321 1008
rect 3334 961 3337 968
rect 3334 958 3345 961
rect 3342 952 3345 958
rect 3358 952 3361 1058
rect 3390 1052 3393 1058
rect 3454 1052 3457 1058
rect 3406 1042 3409 1048
rect 3374 968 3382 971
rect 3366 962 3369 968
rect 3322 878 3326 881
rect 3322 868 3326 871
rect 3334 862 3337 948
rect 3366 942 3369 948
rect 3346 938 3350 941
rect 3374 892 3377 968
rect 3382 942 3385 958
rect 3390 952 3393 1018
rect 3398 962 3401 1028
rect 3486 1022 3489 1068
rect 3494 1052 3497 1108
rect 3502 1062 3505 1068
rect 3502 1042 3505 1048
rect 3408 1003 3410 1007
rect 3414 1003 3417 1007
rect 3421 1003 3424 1007
rect 3402 948 3406 951
rect 3422 932 3425 978
rect 3494 972 3497 978
rect 3502 972 3505 1038
rect 3510 992 3513 1068
rect 3478 968 3486 971
rect 3470 962 3473 968
rect 3446 932 3449 938
rect 3470 912 3473 918
rect 3406 882 3409 888
rect 3378 878 3382 881
rect 3478 872 3481 968
rect 3506 958 3510 961
rect 3490 948 3494 951
rect 3502 872 3505 948
rect 3518 942 3521 1108
rect 3542 1102 3545 1138
rect 3550 1092 3553 1168
rect 3558 1152 3561 1278
rect 3586 1268 3590 1271
rect 3566 1262 3569 1268
rect 3582 1252 3585 1258
rect 3606 1252 3609 1268
rect 3662 1262 3665 1268
rect 3670 1262 3673 1308
rect 3678 1302 3681 1338
rect 3678 1272 3681 1288
rect 3566 1162 3569 1168
rect 3566 1082 3569 1148
rect 3574 1142 3577 1238
rect 3606 1191 3609 1248
rect 3618 1238 3622 1241
rect 3630 1231 3633 1258
rect 3638 1252 3641 1258
rect 3678 1252 3681 1258
rect 3650 1248 3657 1251
rect 3598 1188 3609 1191
rect 3614 1228 3633 1231
rect 3614 1192 3617 1228
rect 3626 1218 3630 1221
rect 3586 1158 3590 1161
rect 3554 1078 3558 1081
rect 3562 1068 3566 1071
rect 3534 1062 3537 1068
rect 3582 1061 3585 1158
rect 3598 1112 3601 1188
rect 3606 1172 3609 1178
rect 3618 1158 3622 1161
rect 3614 1142 3617 1148
rect 3630 1142 3633 1208
rect 3594 1088 3598 1091
rect 3578 1058 3585 1061
rect 3526 1002 3529 1048
rect 3550 992 3553 1058
rect 3590 1052 3593 1078
rect 3602 1068 3606 1071
rect 3618 1068 3622 1071
rect 3630 1062 3633 1128
rect 3614 1042 3617 1048
rect 3622 1042 3625 1058
rect 3582 972 3585 978
rect 3590 972 3593 1038
rect 3614 992 3617 1028
rect 3630 1022 3633 1028
rect 3606 972 3609 978
rect 3526 942 3529 948
rect 3510 922 3513 928
rect 3518 892 3521 918
rect 3526 882 3529 898
rect 3346 868 3350 871
rect 3402 868 3406 871
rect 3458 868 3462 871
rect 3510 862 3513 868
rect 3346 858 3350 861
rect 3458 858 3462 861
rect 3318 842 3321 858
rect 3358 852 3361 858
rect 3378 848 3382 851
rect 3342 842 3345 848
rect 3310 838 3318 841
rect 3282 748 3286 751
rect 3262 742 3265 748
rect 3206 732 3209 738
rect 3246 732 3249 738
rect 3278 732 3281 748
rect 3226 728 3230 731
rect 3174 722 3177 728
rect 3162 718 3166 721
rect 3214 702 3217 718
rect 3158 672 3161 678
rect 3214 672 3217 678
rect 3254 672 3257 708
rect 3262 682 3265 688
rect 3162 658 3166 661
rect 3202 658 3206 661
rect 3222 652 3225 658
rect 3158 562 3161 608
rect 3182 602 3185 618
rect 3190 612 3193 648
rect 3238 622 3241 658
rect 3174 572 3177 578
rect 3158 552 3161 558
rect 3170 548 3174 551
rect 3182 542 3185 558
rect 3206 551 3209 618
rect 3238 572 3241 618
rect 3254 582 3257 668
rect 3270 661 3273 718
rect 3286 662 3289 678
rect 3294 672 3297 818
rect 3330 748 3334 751
rect 3350 751 3353 838
rect 3374 762 3377 848
rect 3398 842 3401 858
rect 3470 852 3473 858
rect 3454 842 3457 848
rect 3408 803 3410 807
rect 3414 803 3417 807
rect 3421 803 3424 807
rect 3434 788 3438 791
rect 3446 762 3449 838
rect 3462 762 3465 768
rect 3382 752 3385 758
rect 3478 752 3481 858
rect 3518 852 3521 868
rect 3486 842 3489 848
rect 3486 752 3489 758
rect 3346 748 3353 751
rect 3394 748 3398 751
rect 3306 738 3310 741
rect 3330 728 3334 731
rect 3302 722 3305 728
rect 3310 692 3313 728
rect 3318 722 3321 728
rect 3310 662 3313 668
rect 3270 658 3281 661
rect 3270 642 3273 648
rect 3214 562 3217 568
rect 3202 548 3209 551
rect 3214 542 3217 548
rect 3222 542 3225 548
rect 3238 541 3241 568
rect 3234 538 3241 541
rect 3190 532 3193 538
rect 3190 472 3193 528
rect 3230 502 3233 538
rect 3238 482 3241 518
rect 3254 481 3257 558
rect 3270 532 3273 548
rect 3278 542 3281 658
rect 3326 652 3329 678
rect 3342 671 3345 748
rect 3358 742 3361 748
rect 3474 738 3478 741
rect 3350 731 3353 738
rect 3350 728 3361 731
rect 3358 692 3361 728
rect 3374 692 3377 728
rect 3382 722 3385 728
rect 3398 692 3401 738
rect 3422 732 3425 738
rect 3450 728 3454 731
rect 3462 692 3465 718
rect 3494 692 3497 848
rect 3518 792 3521 818
rect 3542 792 3545 968
rect 3550 952 3553 958
rect 3558 932 3561 958
rect 3574 922 3577 968
rect 3590 962 3593 968
rect 3582 912 3585 948
rect 3590 892 3593 918
rect 3558 872 3561 888
rect 3562 858 3566 861
rect 3574 852 3577 858
rect 3558 842 3561 848
rect 3582 792 3585 878
rect 3590 842 3593 848
rect 3602 828 3606 831
rect 3614 792 3617 948
rect 3622 932 3625 958
rect 3638 941 3641 1228
rect 3646 1142 3649 1158
rect 3646 1132 3649 1138
rect 3646 1062 3649 1118
rect 3646 1042 3649 1048
rect 3654 1022 3657 1248
rect 3662 1042 3665 1048
rect 3670 992 3673 1228
rect 3686 1152 3689 1478
rect 3702 1462 3705 1468
rect 3718 1462 3721 1468
rect 3694 1432 3697 1448
rect 3702 1372 3705 1378
rect 3694 1342 3697 1368
rect 3710 1362 3713 1418
rect 3718 1392 3721 1438
rect 3726 1422 3729 1558
rect 3746 1548 3750 1551
rect 3758 1541 3761 1628
rect 3750 1538 3761 1541
rect 3750 1442 3753 1538
rect 3758 1452 3761 1458
rect 3742 1422 3745 1428
rect 3726 1372 3729 1378
rect 3734 1352 3737 1408
rect 3742 1362 3745 1368
rect 3758 1352 3761 1398
rect 3766 1392 3769 1648
rect 3774 1372 3777 1638
rect 3770 1358 3774 1361
rect 3706 1348 3710 1351
rect 3770 1348 3774 1351
rect 3750 1332 3753 1338
rect 3694 1242 3697 1318
rect 3706 1278 3710 1281
rect 3718 1261 3721 1278
rect 3726 1272 3729 1298
rect 3742 1272 3745 1278
rect 3758 1272 3761 1288
rect 3706 1258 3721 1261
rect 3730 1258 3734 1261
rect 3738 1248 3742 1251
rect 3750 1192 3753 1248
rect 3758 1202 3761 1258
rect 3822 1222 3825 1838
rect 3726 1172 3729 1178
rect 3754 1168 3758 1171
rect 3742 1152 3745 1158
rect 3678 1072 3681 1148
rect 3686 1102 3689 1148
rect 3726 1142 3729 1148
rect 3686 1072 3689 1088
rect 3702 1082 3705 1118
rect 3710 1092 3713 1138
rect 3742 1092 3745 1138
rect 3678 1062 3681 1068
rect 3694 1002 3697 1058
rect 3662 972 3665 988
rect 3634 938 3641 941
rect 3646 962 3649 968
rect 3674 958 3678 961
rect 3622 832 3625 928
rect 3638 882 3641 918
rect 3634 868 3638 871
rect 3646 861 3649 958
rect 3686 952 3689 958
rect 3670 932 3673 948
rect 3686 912 3689 938
rect 3694 912 3697 998
rect 3710 962 3713 1058
rect 3718 1032 3721 1068
rect 3726 952 3729 1058
rect 3726 942 3729 948
rect 3642 858 3649 861
rect 3630 852 3633 858
rect 3502 762 3505 768
rect 3526 758 3534 761
rect 3514 748 3518 751
rect 3502 732 3505 738
rect 3510 702 3513 738
rect 3362 678 3366 681
rect 3426 678 3430 681
rect 3338 668 3345 671
rect 3334 662 3337 668
rect 3378 658 3382 661
rect 3286 642 3289 648
rect 3342 632 3345 658
rect 3286 542 3289 598
rect 3306 558 3310 561
rect 3294 522 3297 548
rect 3326 542 3329 618
rect 3390 612 3393 678
rect 3402 658 3406 661
rect 3434 658 3438 661
rect 3408 603 3410 607
rect 3414 603 3417 607
rect 3421 603 3424 607
rect 3334 542 3337 568
rect 3342 552 3345 598
rect 3382 562 3385 578
rect 3354 548 3358 551
rect 3346 538 3350 541
rect 3262 492 3265 518
rect 3326 482 3329 518
rect 3254 478 3265 481
rect 3262 472 3265 478
rect 3302 472 3305 478
rect 3266 468 3270 471
rect 3094 362 3097 458
rect 3106 388 3110 391
rect 3150 372 3153 458
rect 3182 431 3185 450
rect 3162 358 3166 361
rect 3054 212 3057 268
rect 3078 262 3081 338
rect 3110 312 3113 318
rect 3110 292 3113 308
rect 3098 248 3102 251
rect 3126 232 3129 348
rect 3134 332 3137 338
rect 3150 332 3153 358
rect 3162 338 3166 341
rect 3174 332 3177 348
rect 3190 342 3193 468
rect 3226 458 3230 461
rect 3222 402 3225 448
rect 3214 362 3217 368
rect 3198 342 3201 348
rect 3226 338 3230 341
rect 3182 332 3185 338
rect 3142 252 3145 318
rect 3150 302 3153 328
rect 3190 272 3193 278
rect 3206 272 3209 278
rect 3150 262 3153 268
rect 3062 202 3065 218
rect 3066 188 3070 191
rect 3078 162 3081 218
rect 3010 158 3014 161
rect 2994 148 2998 151
rect 3010 148 3014 151
rect 3038 142 3041 158
rect 3046 142 3049 148
rect 2994 138 2998 141
rect 3026 138 3030 141
rect 2904 103 2906 107
rect 2910 103 2913 107
rect 2917 103 2920 107
rect 2950 62 2953 118
rect 3006 82 3009 128
rect 3022 122 3025 128
rect 3086 92 3089 208
rect 3094 92 3097 118
rect 3102 82 3105 198
rect 3190 152 3193 258
rect 3206 162 3209 188
rect 3238 182 3241 458
rect 3254 412 3257 468
rect 3350 462 3353 498
rect 3358 472 3361 518
rect 3374 472 3377 518
rect 3382 492 3385 558
rect 3446 552 3449 658
rect 3454 632 3457 668
rect 3478 662 3481 688
rect 3486 672 3489 688
rect 3506 678 3510 681
rect 3518 672 3521 748
rect 3526 692 3529 758
rect 3542 692 3545 778
rect 3622 772 3625 788
rect 3550 762 3553 768
rect 3590 758 3598 761
rect 3534 672 3537 678
rect 3558 672 3561 748
rect 3566 712 3569 758
rect 3582 752 3585 758
rect 3574 722 3577 738
rect 3474 648 3478 651
rect 3454 592 3457 608
rect 3442 548 3446 551
rect 3398 502 3401 548
rect 3406 522 3409 538
rect 3446 532 3449 538
rect 3462 532 3465 618
rect 3510 612 3513 658
rect 3518 652 3521 668
rect 3542 661 3545 668
rect 3574 662 3577 698
rect 3582 672 3585 748
rect 3590 692 3593 758
rect 3606 712 3609 758
rect 3614 732 3617 748
rect 3606 682 3609 688
rect 3598 672 3601 678
rect 3534 658 3545 661
rect 3554 658 3558 661
rect 3534 592 3537 658
rect 3566 652 3569 658
rect 3574 652 3577 658
rect 3582 652 3585 668
rect 3566 572 3569 648
rect 3602 618 3606 621
rect 3614 592 3617 708
rect 3630 702 3633 778
rect 3638 742 3641 808
rect 3646 792 3649 858
rect 3654 852 3657 878
rect 3690 868 3694 871
rect 3662 862 3665 868
rect 3702 862 3705 868
rect 3670 822 3673 858
rect 3670 782 3673 818
rect 3686 802 3689 858
rect 3702 842 3705 858
rect 3710 832 3713 908
rect 3718 892 3721 928
rect 3722 868 3726 871
rect 3734 861 3737 1078
rect 3758 962 3761 1018
rect 3766 952 3769 1148
rect 3774 1122 3777 1158
rect 3774 1062 3777 1068
rect 3774 952 3777 958
rect 3750 932 3753 938
rect 3726 858 3737 861
rect 3746 858 3750 861
rect 3654 762 3657 778
rect 3686 772 3689 788
rect 3662 768 3670 771
rect 3654 742 3657 748
rect 3662 731 3665 768
rect 3686 762 3689 768
rect 3674 748 3678 751
rect 3686 741 3689 748
rect 3682 738 3689 741
rect 3654 728 3665 731
rect 3690 728 3694 731
rect 3630 672 3633 698
rect 3566 562 3569 568
rect 3598 562 3601 568
rect 3610 558 3614 561
rect 3470 552 3473 558
rect 3490 548 3494 551
rect 3514 548 3518 551
rect 3554 548 3558 551
rect 3570 548 3574 551
rect 3610 548 3614 551
rect 3510 532 3513 538
rect 3518 532 3521 538
rect 3426 528 3430 531
rect 3482 528 3486 531
rect 3494 512 3497 528
rect 3534 522 3537 548
rect 3582 542 3585 548
rect 3598 542 3601 548
rect 3566 538 3574 541
rect 3542 532 3545 538
rect 3566 492 3569 538
rect 3538 488 3542 491
rect 3446 472 3449 478
rect 3462 472 3465 478
rect 3274 458 3278 461
rect 3290 448 3294 451
rect 3246 272 3249 318
rect 3254 312 3257 358
rect 3270 352 3273 438
rect 3302 362 3305 378
rect 3270 302 3273 348
rect 3278 342 3281 348
rect 3278 302 3281 318
rect 3286 312 3289 338
rect 3302 332 3305 338
rect 3294 322 3297 328
rect 3310 312 3313 418
rect 3334 412 3337 448
rect 3350 442 3353 458
rect 3338 408 3345 411
rect 3330 358 3334 361
rect 3270 282 3273 298
rect 3278 272 3281 298
rect 3318 292 3321 348
rect 3330 338 3334 341
rect 3342 282 3345 408
rect 3350 362 3353 368
rect 3358 352 3361 468
rect 3366 362 3369 468
rect 3382 352 3385 418
rect 3390 352 3393 448
rect 3398 422 3401 448
rect 3408 403 3410 407
rect 3414 403 3417 407
rect 3421 403 3424 407
rect 3446 352 3449 438
rect 3502 411 3505 458
rect 3494 408 3505 411
rect 3466 358 3470 361
rect 3486 352 3489 368
rect 3474 348 3478 351
rect 3350 332 3353 348
rect 3382 342 3385 348
rect 3390 342 3393 348
rect 3438 342 3441 348
rect 3426 338 3430 341
rect 3474 338 3478 341
rect 3374 332 3377 338
rect 3406 302 3409 338
rect 3418 328 3422 331
rect 3446 282 3449 288
rect 3330 278 3334 281
rect 3462 272 3465 308
rect 3318 262 3321 268
rect 3282 258 3286 261
rect 3254 222 3257 248
rect 3302 242 3305 248
rect 3282 218 3286 221
rect 3302 192 3305 228
rect 3310 202 3313 258
rect 3326 252 3329 258
rect 3158 142 3161 148
rect 3142 132 3145 138
rect 3110 92 3113 98
rect 3126 92 3129 108
rect 3146 88 3150 91
rect 3138 78 3142 81
rect 2990 72 2993 78
rect 3190 72 3193 148
rect 3226 138 3230 141
rect 3290 138 3294 141
rect 3230 82 3233 128
rect 3246 72 3249 78
rect 3046 62 3049 68
rect 3190 62 3193 68
rect 3302 62 3305 138
rect 3310 122 3313 138
rect 3334 92 3337 268
rect 3494 262 3497 408
rect 3510 392 3513 418
rect 3534 392 3537 478
rect 3558 422 3561 478
rect 3574 462 3577 518
rect 3622 501 3625 568
rect 3630 512 3633 658
rect 3638 632 3641 668
rect 3646 592 3649 718
rect 3654 692 3657 728
rect 3662 662 3665 668
rect 3682 648 3686 651
rect 3654 612 3657 648
rect 3678 592 3681 628
rect 3694 622 3697 668
rect 3702 642 3705 828
rect 3726 792 3729 858
rect 3726 772 3729 778
rect 3710 761 3713 768
rect 3734 761 3737 828
rect 3754 768 3758 771
rect 3710 758 3721 761
rect 3718 752 3721 758
rect 3734 758 3742 761
rect 3770 758 3774 761
rect 3710 742 3713 748
rect 3710 692 3713 718
rect 3718 712 3721 738
rect 3710 672 3713 678
rect 3726 672 3729 678
rect 3642 558 3646 561
rect 3646 542 3649 548
rect 3622 498 3633 501
rect 3630 492 3633 498
rect 3582 482 3585 488
rect 3598 472 3601 478
rect 3654 472 3657 568
rect 3670 502 3673 528
rect 3670 482 3673 488
rect 3594 458 3598 461
rect 3502 352 3505 358
rect 3518 342 3521 358
rect 3574 342 3577 458
rect 3502 282 3505 318
rect 3408 203 3410 207
rect 3414 203 3417 207
rect 3421 203 3424 207
rect 3366 142 3369 148
rect 3406 142 3409 188
rect 3422 142 3425 148
rect 3406 132 3409 138
rect 3354 68 3358 71
rect 3334 62 3337 68
rect 3390 62 3393 68
rect 2226 58 2230 61
rect 2562 58 2566 61
rect 2738 58 2742 61
rect 2850 58 2854 61
rect 2906 58 2910 61
rect 3122 58 3126 61
rect 1870 31 1873 50
rect 1926 -18 1929 8
rect 1998 -18 2001 28
rect 2046 22 2049 50
rect 2246 22 2249 50
rect 2410 48 2414 51
rect 3366 52 3369 58
rect 3398 52 3401 98
rect 3454 92 3457 208
rect 3462 152 3465 258
rect 3494 252 3497 258
rect 3470 162 3473 188
rect 3502 92 3505 268
rect 3510 222 3513 248
rect 3518 192 3521 318
rect 3534 222 3537 268
rect 3534 152 3537 208
rect 3430 82 3433 88
rect 3446 62 3449 88
rect 3470 62 3473 68
rect 3486 62 3489 78
rect 3526 62 3529 68
rect 3542 62 3545 178
rect 3554 168 3558 171
rect 3566 162 3569 168
rect 3554 148 3558 151
rect 3574 122 3577 338
rect 3582 192 3585 438
rect 3606 432 3609 468
rect 3614 462 3617 468
rect 3626 448 3630 451
rect 3638 442 3641 468
rect 3646 462 3649 468
rect 3658 448 3662 451
rect 3590 292 3593 338
rect 3598 322 3601 328
rect 3590 192 3593 218
rect 3598 152 3601 158
rect 3550 72 3553 118
rect 3574 72 3577 118
rect 3598 92 3601 148
rect 3606 142 3609 408
rect 3614 392 3617 438
rect 3630 392 3633 428
rect 3678 392 3681 558
rect 3686 552 3689 608
rect 3690 548 3694 551
rect 3694 512 3697 528
rect 3702 512 3705 598
rect 3710 522 3713 548
rect 3718 542 3721 548
rect 3718 522 3721 528
rect 3686 462 3689 468
rect 3702 462 3705 488
rect 3710 472 3713 518
rect 3718 492 3721 508
rect 3726 482 3729 648
rect 3734 582 3737 758
rect 3762 748 3766 751
rect 3750 692 3753 718
rect 3758 672 3761 678
rect 3742 662 3745 668
rect 3750 652 3753 658
rect 3762 648 3766 651
rect 3750 592 3753 638
rect 3734 561 3737 568
rect 3766 562 3769 568
rect 3734 558 3745 561
rect 3742 552 3745 558
rect 3734 492 3737 548
rect 3742 532 3745 538
rect 3742 492 3745 498
rect 3774 481 3777 668
rect 3770 478 3777 481
rect 3726 471 3729 478
rect 3718 468 3729 471
rect 3698 458 3702 461
rect 3718 432 3721 468
rect 3734 462 3737 468
rect 3726 392 3729 458
rect 3634 358 3638 361
rect 3614 292 3617 358
rect 3646 352 3649 368
rect 3654 352 3657 358
rect 3662 352 3665 358
rect 3622 342 3625 348
rect 3622 322 3625 328
rect 3606 82 3609 108
rect 3614 92 3617 258
rect 3626 148 3630 151
rect 3638 92 3641 328
rect 3646 322 3649 348
rect 3646 192 3649 298
rect 3630 82 3633 88
rect 3586 68 3590 71
rect 3654 62 3657 348
rect 3758 342 3761 348
rect 3666 338 3670 341
rect 3706 338 3710 341
rect 3694 282 3697 288
rect 3710 272 3713 278
rect 3710 252 3713 258
rect 3742 231 3745 250
rect 3718 192 3721 218
rect 3758 212 3761 318
rect 3766 232 3769 478
rect 3742 192 3745 198
rect 3714 168 3718 171
rect 3662 152 3665 158
rect 3718 152 3721 158
rect 3674 148 3678 151
rect 3674 138 3678 141
rect 3726 141 3729 158
rect 3758 152 3761 208
rect 3718 138 3729 141
rect 3698 128 3702 131
rect 3662 92 3665 128
rect 3686 92 3689 118
rect 3694 81 3697 108
rect 3718 102 3721 138
rect 3718 92 3721 98
rect 3686 78 3697 81
rect 3722 78 3726 81
rect 3686 72 3689 78
rect 3698 68 3702 71
rect 3678 62 3681 68
rect 3618 58 3622 61
rect 3690 58 3694 61
rect 3478 52 3481 58
rect 3646 52 3649 58
rect 3710 52 3713 58
rect 3726 52 3729 58
rect 3734 52 3737 88
rect 3758 72 3761 78
rect 2542 31 2545 50
rect 3354 48 3358 51
rect 2734 22 2737 48
rect 2942 22 2945 48
rect 3294 22 3297 48
rect 3330 38 3334 41
rect 3342 32 3345 48
rect 3750 42 3753 58
rect 3378 38 3382 41
rect 3458 38 3462 41
rect 3390 32 3393 38
rect 3590 32 3593 38
rect 2094 -18 2097 8
rect 2384 3 2386 7
rect 2390 3 2393 7
rect 2397 3 2400 7
rect 2494 -18 2497 8
rect 3408 3 3410 7
rect 3414 3 3417 7
rect 3421 3 3424 7
rect 1862 -22 1866 -18
rect 1926 -22 1930 -18
rect 1998 -22 2002 -18
rect 2094 -22 2098 -18
rect 2494 -22 2498 -18
<< m3contact >>
rect 30 3538 34 3542
rect 62 3538 66 3542
rect 86 3538 90 3542
rect 102 3538 106 3542
rect 174 3538 178 3542
rect 6 3468 10 3472
rect 6 3448 10 3452
rect 166 3478 170 3482
rect 86 3428 90 3432
rect 134 3428 138 3432
rect 346 3603 350 3607
rect 353 3603 357 3607
rect 430 3598 434 3602
rect 886 3598 890 3602
rect 318 3548 322 3552
rect 374 3548 378 3552
rect 518 3548 522 3552
rect 606 3548 610 3552
rect 726 3548 730 3552
rect 238 3528 242 3532
rect 198 3448 202 3452
rect 174 3408 178 3412
rect 22 3398 26 3402
rect 182 3388 186 3392
rect 6 3378 10 3382
rect 286 3518 290 3522
rect 318 3468 322 3472
rect 334 3458 338 3462
rect 294 3408 298 3412
rect 346 3403 350 3407
rect 353 3403 357 3407
rect 326 3398 330 3402
rect 446 3518 450 3522
rect 422 3508 426 3512
rect 438 3448 442 3452
rect 454 3398 458 3402
rect 286 3388 290 3392
rect 318 3388 322 3392
rect 358 3388 362 3392
rect 382 3388 386 3392
rect 246 3368 250 3372
rect 30 3358 34 3362
rect 22 3348 26 3352
rect 246 3348 250 3352
rect 6 3248 10 3252
rect 14 3138 18 3142
rect 6 3048 10 3052
rect 6 2948 10 2952
rect 54 3338 58 3342
rect 70 3338 74 3342
rect 62 3328 66 3332
rect 174 3318 178 3322
rect 350 3358 354 3362
rect 318 3348 322 3352
rect 310 3338 314 3342
rect 254 3328 258 3332
rect 270 3328 274 3332
rect 262 3318 266 3322
rect 134 3258 138 3262
rect 118 3248 122 3252
rect 134 3248 138 3252
rect 22 3078 26 3082
rect 46 3078 50 3082
rect 22 3048 26 3052
rect 174 3308 178 3312
rect 206 3308 210 3312
rect 278 3308 282 3312
rect 222 3298 226 3302
rect 286 3298 290 3302
rect 318 3298 322 3302
rect 206 3238 210 3242
rect 406 3378 410 3382
rect 454 3368 458 3372
rect 366 3348 370 3352
rect 422 3348 426 3352
rect 398 3338 402 3342
rect 390 3328 394 3332
rect 366 3298 370 3302
rect 374 3298 378 3302
rect 414 3318 418 3322
rect 406 3288 410 3292
rect 366 3278 370 3282
rect 318 3248 322 3252
rect 302 3228 306 3232
rect 206 3218 210 3222
rect 446 3328 450 3332
rect 446 3258 450 3262
rect 438 3248 442 3252
rect 422 3238 426 3242
rect 346 3203 350 3207
rect 353 3203 357 3207
rect 214 3158 218 3162
rect 166 3128 170 3132
rect 134 3058 138 3062
rect 86 3008 90 3012
rect 118 3008 122 3012
rect 454 3208 458 3212
rect 278 3148 282 3152
rect 294 3148 298 3152
rect 366 3148 370 3152
rect 406 3148 410 3152
rect 230 3118 234 3122
rect 254 3098 258 3102
rect 206 3078 210 3082
rect 230 3078 234 3082
rect 214 3068 218 3072
rect 238 3068 242 3072
rect 230 3058 234 3062
rect 246 3048 250 3052
rect 230 3038 234 3042
rect 78 2938 82 2942
rect 94 2938 98 2942
rect 166 2938 170 2942
rect 238 2938 242 2942
rect 22 2928 26 2932
rect 238 2928 242 2932
rect 30 2908 34 2912
rect 70 2908 74 2912
rect 30 2888 34 2892
rect 54 2878 58 2882
rect 14 2868 18 2872
rect 6 2848 10 2852
rect 6 2748 10 2752
rect 6 2668 10 2672
rect 6 2558 10 2562
rect 6 2488 10 2492
rect 6 2468 10 2472
rect 6 2448 10 2452
rect 6 2348 10 2352
rect 30 2858 34 2862
rect 54 2858 58 2862
rect 46 2848 50 2852
rect 62 2838 66 2842
rect 70 2818 74 2822
rect 54 2798 58 2802
rect 94 2888 98 2892
rect 118 2878 122 2882
rect 118 2858 122 2862
rect 110 2848 114 2852
rect 134 2848 138 2852
rect 86 2808 90 2812
rect 206 2868 210 2872
rect 230 2868 234 2872
rect 422 3118 426 3122
rect 310 3098 314 3102
rect 342 3058 346 3062
rect 446 3068 450 3072
rect 454 3048 458 3052
rect 358 3028 362 3032
rect 346 3003 350 3007
rect 353 3003 357 3007
rect 334 2938 338 2942
rect 310 2928 314 2932
rect 414 2938 418 2942
rect 342 2898 346 2902
rect 214 2858 218 2862
rect 254 2848 258 2852
rect 158 2828 162 2832
rect 230 2828 234 2832
rect 374 2858 378 2862
rect 166 2818 170 2822
rect 94 2798 98 2802
rect 142 2798 146 2802
rect 134 2748 138 2752
rect 78 2708 82 2712
rect 70 2668 74 2672
rect 214 2708 218 2712
rect 318 2828 322 2832
rect 294 2808 298 2812
rect 346 2803 350 2807
rect 353 2803 357 2807
rect 342 2758 346 2762
rect 310 2748 314 2752
rect 374 2738 378 2742
rect 294 2728 298 2732
rect 318 2708 322 2712
rect 214 2678 218 2682
rect 534 3488 538 3492
rect 662 3528 666 3532
rect 902 3528 906 3532
rect 702 3518 706 3522
rect 886 3518 890 3522
rect 646 3488 650 3492
rect 850 3503 854 3507
rect 857 3503 861 3507
rect 606 3458 610 3462
rect 630 3458 634 3462
rect 550 3408 554 3412
rect 646 3448 650 3452
rect 598 3408 602 3412
rect 518 3318 522 3322
rect 534 3318 538 3322
rect 550 3308 554 3312
rect 470 3298 474 3302
rect 518 3288 522 3292
rect 478 3278 482 3282
rect 510 3268 514 3272
rect 670 3408 674 3412
rect 654 3398 658 3402
rect 606 3338 610 3342
rect 614 3328 618 3332
rect 630 3308 634 3312
rect 622 3298 626 3302
rect 646 3298 650 3302
rect 662 3318 666 3322
rect 1070 3598 1074 3602
rect 1078 3568 1082 3572
rect 958 3528 962 3532
rect 894 3458 898 3462
rect 886 3378 890 3382
rect 878 3368 882 3372
rect 870 3358 874 3362
rect 782 3338 786 3342
rect 830 3338 834 3342
rect 782 3318 786 3322
rect 694 3308 698 3312
rect 702 3308 706 3312
rect 774 3308 778 3312
rect 686 3298 690 3302
rect 766 3298 770 3302
rect 558 3268 562 3272
rect 606 3268 610 3272
rect 678 3268 682 3272
rect 686 3268 690 3272
rect 702 3268 706 3272
rect 534 3248 538 3252
rect 566 3248 570 3252
rect 478 3238 482 3242
rect 486 3208 490 3212
rect 486 3068 490 3072
rect 462 2898 466 2902
rect 502 3018 506 3022
rect 526 3238 530 3242
rect 622 3258 626 3262
rect 598 3248 602 3252
rect 630 3218 634 3222
rect 582 3178 586 3182
rect 518 3148 522 3152
rect 526 3148 530 3152
rect 582 3148 586 3152
rect 526 3138 530 3142
rect 518 3048 522 3052
rect 494 2998 498 3002
rect 598 3118 602 3122
rect 582 3088 586 3092
rect 566 3078 570 3082
rect 622 3028 626 3032
rect 678 3198 682 3202
rect 710 3258 714 3262
rect 782 3278 786 3282
rect 846 3328 850 3332
rect 850 3303 854 3307
rect 857 3303 861 3307
rect 878 3348 882 3352
rect 886 3308 890 3312
rect 870 3298 874 3302
rect 806 3268 810 3272
rect 814 3258 818 3262
rect 758 3248 762 3252
rect 718 3238 722 3242
rect 718 3218 722 3222
rect 694 3198 698 3202
rect 750 3168 754 3172
rect 702 3148 706 3152
rect 718 3138 722 3142
rect 774 3178 778 3182
rect 742 3158 746 3162
rect 766 3158 770 3162
rect 710 3128 714 3132
rect 734 3128 738 3132
rect 670 3058 674 3062
rect 670 3038 674 3042
rect 622 3018 626 3022
rect 598 2988 602 2992
rect 574 2978 578 2982
rect 542 2968 546 2972
rect 518 2958 522 2962
rect 558 2958 562 2962
rect 550 2948 554 2952
rect 502 2918 506 2922
rect 534 2928 538 2932
rect 526 2908 530 2912
rect 574 2948 578 2952
rect 574 2918 578 2922
rect 566 2888 570 2892
rect 478 2868 482 2872
rect 422 2858 426 2862
rect 454 2858 458 2862
rect 510 2858 514 2862
rect 414 2808 418 2812
rect 422 2718 426 2722
rect 398 2708 402 2712
rect 366 2688 370 2692
rect 462 2778 466 2782
rect 550 2808 554 2812
rect 542 2768 546 2772
rect 478 2738 482 2742
rect 526 2738 530 2742
rect 422 2678 426 2682
rect 430 2678 434 2682
rect 406 2668 410 2672
rect 478 2708 482 2712
rect 518 2708 522 2712
rect 462 2688 466 2692
rect 318 2658 322 2662
rect 342 2658 346 2662
rect 358 2658 362 2662
rect 382 2658 386 2662
rect 398 2658 402 2662
rect 118 2578 122 2582
rect 366 2648 370 2652
rect 382 2648 386 2652
rect 366 2608 370 2612
rect 346 2603 350 2607
rect 353 2603 357 2607
rect 414 2648 418 2652
rect 390 2588 394 2592
rect 134 2548 138 2552
rect 366 2548 370 2552
rect 182 2538 186 2542
rect 254 2538 258 2542
rect 294 2538 298 2542
rect 78 2528 82 2532
rect 118 2518 122 2522
rect 174 2518 178 2522
rect 222 2518 226 2522
rect 134 2508 138 2512
rect 62 2488 66 2492
rect 30 2478 34 2482
rect 54 2478 58 2482
rect 102 2478 106 2482
rect 86 2468 90 2472
rect 30 2458 34 2462
rect 54 2458 58 2462
rect 46 2448 50 2452
rect 30 2378 34 2382
rect 86 2448 90 2452
rect 62 2438 66 2442
rect 54 2308 58 2312
rect 62 2308 66 2312
rect 22 2278 26 2282
rect 14 2268 18 2272
rect 38 2268 42 2272
rect 54 2268 58 2272
rect 6 2248 10 2252
rect 22 2248 26 2252
rect 46 2188 50 2192
rect 6 2148 10 2152
rect 6 2078 10 2082
rect 30 2048 34 2052
rect 22 2038 26 2042
rect 54 2068 58 2072
rect 190 2458 194 2462
rect 174 2418 178 2422
rect 198 2418 202 2422
rect 110 2308 114 2312
rect 102 2268 106 2272
rect 110 2268 114 2272
rect 158 2318 162 2322
rect 294 2448 298 2452
rect 414 2528 418 2532
rect 366 2488 370 2492
rect 382 2488 386 2492
rect 310 2428 314 2432
rect 346 2403 350 2407
rect 353 2403 357 2407
rect 294 2368 298 2372
rect 214 2348 218 2352
rect 238 2348 242 2352
rect 358 2348 362 2352
rect 454 2658 458 2662
rect 510 2658 514 2662
rect 542 2658 546 2662
rect 502 2648 506 2652
rect 446 2638 450 2642
rect 478 2638 482 2642
rect 486 2638 490 2642
rect 502 2638 506 2642
rect 446 2548 450 2552
rect 502 2548 506 2552
rect 438 2468 442 2472
rect 478 2508 482 2512
rect 462 2498 466 2502
rect 438 2458 442 2462
rect 446 2458 450 2462
rect 454 2448 458 2452
rect 470 2448 474 2452
rect 438 2438 442 2442
rect 382 2348 386 2352
rect 310 2308 314 2312
rect 326 2308 330 2312
rect 366 2308 370 2312
rect 326 2288 330 2292
rect 198 2278 202 2282
rect 342 2278 346 2282
rect 206 2268 210 2272
rect 254 2268 258 2272
rect 94 2258 98 2262
rect 134 2258 138 2262
rect 142 2258 146 2262
rect 238 2258 242 2262
rect 118 2248 122 2252
rect 134 2248 138 2252
rect 86 2208 90 2212
rect 118 2208 122 2212
rect 134 2148 138 2152
rect 118 2118 122 2122
rect 78 2068 82 2072
rect 206 2128 210 2132
rect 446 2388 450 2392
rect 454 2358 458 2362
rect 606 2948 610 2952
rect 598 2938 602 2942
rect 598 2878 602 2882
rect 694 2998 698 3002
rect 742 3118 746 3122
rect 734 3068 738 3072
rect 742 3058 746 3062
rect 734 3048 738 3052
rect 798 3168 802 3172
rect 798 3158 802 3162
rect 766 3128 770 3132
rect 774 3128 778 3132
rect 782 3108 786 3112
rect 774 3098 778 3102
rect 774 3078 778 3082
rect 830 3178 834 3182
rect 878 3168 882 3172
rect 870 3158 874 3162
rect 878 3158 882 3162
rect 838 3148 842 3152
rect 846 3138 850 3142
rect 822 3118 826 3122
rect 850 3103 854 3107
rect 857 3103 861 3107
rect 798 3078 802 3082
rect 782 3068 786 3072
rect 782 3058 786 3062
rect 710 2988 714 2992
rect 638 2978 642 2982
rect 654 2978 658 2982
rect 678 2978 682 2982
rect 630 2968 634 2972
rect 638 2968 642 2972
rect 694 2968 698 2972
rect 670 2928 674 2932
rect 686 2928 690 2932
rect 638 2918 642 2922
rect 646 2918 650 2922
rect 630 2908 634 2912
rect 654 2888 658 2892
rect 726 2928 730 2932
rect 694 2888 698 2892
rect 702 2888 706 2892
rect 718 2888 722 2892
rect 678 2868 682 2872
rect 598 2848 602 2852
rect 614 2848 618 2852
rect 566 2738 570 2742
rect 582 2688 586 2692
rect 566 2678 570 2682
rect 590 2678 594 2682
rect 646 2788 650 2792
rect 614 2768 618 2772
rect 622 2758 626 2762
rect 614 2748 618 2752
rect 622 2738 626 2742
rect 638 2728 642 2732
rect 630 2698 634 2702
rect 630 2678 634 2682
rect 638 2668 642 2672
rect 574 2658 578 2662
rect 590 2648 594 2652
rect 558 2638 562 2642
rect 574 2638 578 2642
rect 622 2648 626 2652
rect 646 2618 650 2622
rect 662 2798 666 2802
rect 662 2788 666 2792
rect 686 2858 690 2862
rect 678 2838 682 2842
rect 718 2838 722 2842
rect 726 2838 730 2842
rect 766 3038 770 3042
rect 766 3008 770 3012
rect 854 3068 858 3072
rect 846 3058 850 3062
rect 806 3048 810 3052
rect 814 3048 818 3052
rect 830 3048 834 3052
rect 782 2998 786 3002
rect 790 2988 794 2992
rect 758 2978 762 2982
rect 750 2968 754 2972
rect 750 2958 754 2962
rect 766 2938 770 2942
rect 750 2898 754 2902
rect 750 2878 754 2882
rect 774 2878 778 2882
rect 750 2868 754 2872
rect 766 2858 770 2862
rect 774 2858 778 2862
rect 790 2858 794 2862
rect 854 3008 858 3012
rect 862 3008 866 3012
rect 814 2968 818 2972
rect 814 2958 818 2962
rect 830 2948 834 2952
rect 814 2938 818 2942
rect 806 2928 810 2932
rect 814 2898 818 2902
rect 742 2828 746 2832
rect 734 2778 738 2782
rect 718 2768 722 2772
rect 710 2758 714 2762
rect 662 2728 666 2732
rect 670 2708 674 2712
rect 710 2748 714 2752
rect 726 2738 730 2742
rect 742 2738 746 2742
rect 710 2728 714 2732
rect 710 2698 714 2702
rect 726 2668 730 2672
rect 702 2658 706 2662
rect 654 2578 658 2582
rect 670 2578 674 2582
rect 646 2568 650 2572
rect 654 2568 658 2572
rect 718 2648 722 2652
rect 686 2638 690 2642
rect 694 2638 698 2642
rect 782 2828 786 2832
rect 798 2818 802 2822
rect 806 2798 810 2802
rect 806 2788 810 2792
rect 774 2778 778 2782
rect 798 2778 802 2782
rect 758 2768 762 2772
rect 790 2768 794 2772
rect 806 2768 810 2772
rect 774 2758 778 2762
rect 790 2758 794 2762
rect 782 2748 786 2752
rect 774 2688 778 2692
rect 766 2678 770 2682
rect 750 2668 754 2672
rect 742 2648 746 2652
rect 758 2638 762 2642
rect 734 2628 738 2632
rect 782 2678 786 2682
rect 798 2678 802 2682
rect 790 2628 794 2632
rect 822 2868 826 2872
rect 854 2948 858 2952
rect 878 2978 882 2982
rect 870 2958 874 2962
rect 870 2928 874 2932
rect 850 2903 854 2907
rect 857 2903 861 2907
rect 1150 3548 1154 3552
rect 1118 3538 1122 3542
rect 1062 3528 1066 3532
rect 1078 3508 1082 3512
rect 1166 3508 1170 3512
rect 1362 3603 1366 3607
rect 1369 3603 1373 3607
rect 1334 3598 1338 3602
rect 1278 3588 1282 3592
rect 1462 3598 1466 3602
rect 1510 3598 1514 3602
rect 1574 3598 1578 3602
rect 1606 3598 1610 3602
rect 1510 3588 1514 3592
rect 1526 3588 1530 3592
rect 1382 3578 1386 3582
rect 1590 3568 1594 3572
rect 1206 3548 1210 3552
rect 1390 3548 1394 3552
rect 1470 3548 1474 3552
rect 1238 3538 1242 3542
rect 1230 3518 1234 3522
rect 1302 3518 1306 3522
rect 1286 3508 1290 3512
rect 1302 3508 1306 3512
rect 1350 3538 1354 3542
rect 1398 3508 1402 3512
rect 1486 3538 1490 3542
rect 1438 3498 1442 3502
rect 1278 3488 1282 3492
rect 1342 3488 1346 3492
rect 1374 3488 1378 3492
rect 1438 3488 1442 3492
rect 990 3438 994 3442
rect 1054 3428 1058 3432
rect 1062 3418 1066 3422
rect 1054 3408 1058 3412
rect 974 3388 978 3392
rect 998 3378 1002 3382
rect 902 3328 906 3332
rect 950 3358 954 3362
rect 942 3348 946 3352
rect 1046 3348 1050 3352
rect 990 3338 994 3342
rect 1022 3338 1026 3342
rect 1038 3338 1042 3342
rect 926 3308 930 3312
rect 974 3328 978 3332
rect 1222 3468 1226 3472
rect 1246 3468 1250 3472
rect 1270 3468 1274 3472
rect 1302 3468 1306 3472
rect 1214 3458 1218 3462
rect 1086 3388 1090 3392
rect 1222 3448 1226 3452
rect 1158 3428 1162 3432
rect 1190 3428 1194 3432
rect 1758 3598 1762 3602
rect 1662 3548 1666 3552
rect 1574 3528 1578 3532
rect 1630 3528 1634 3532
rect 1750 3528 1754 3532
rect 1902 3598 1906 3602
rect 1974 3598 1978 3602
rect 1790 3588 1794 3592
rect 2386 3603 2390 3607
rect 2393 3603 2397 3607
rect 3410 3603 3414 3607
rect 3417 3603 3421 3607
rect 2230 3598 2234 3602
rect 2406 3598 2410 3602
rect 2078 3588 2082 3592
rect 2430 3588 2434 3592
rect 2902 3588 2906 3592
rect 2942 3588 2946 3592
rect 3262 3588 3266 3592
rect 3342 3588 3346 3592
rect 2062 3568 2066 3572
rect 2022 3558 2026 3562
rect 2262 3568 2266 3572
rect 1990 3548 1994 3552
rect 1814 3538 1818 3542
rect 1798 3528 1802 3532
rect 1854 3528 1858 3532
rect 1742 3478 1746 3482
rect 1614 3468 1618 3472
rect 1262 3458 1266 3462
rect 1286 3458 1290 3462
rect 1310 3458 1314 3462
rect 1422 3458 1426 3462
rect 1478 3458 1482 3462
rect 1526 3458 1530 3462
rect 1542 3458 1546 3462
rect 1262 3438 1266 3442
rect 1246 3398 1250 3402
rect 1230 3368 1234 3372
rect 1110 3348 1114 3352
rect 1126 3348 1130 3352
rect 1070 3318 1074 3322
rect 1190 3328 1194 3332
rect 982 3298 986 3302
rect 1086 3298 1090 3302
rect 942 3268 946 3272
rect 1110 3268 1114 3272
rect 1014 3258 1018 3262
rect 1038 3258 1042 3262
rect 1094 3258 1098 3262
rect 1166 3218 1170 3222
rect 966 3208 970 3212
rect 926 3168 930 3172
rect 1190 3318 1194 3322
rect 1270 3418 1274 3422
rect 1238 3348 1242 3352
rect 1262 3348 1266 3352
rect 1270 3338 1274 3342
rect 1238 3288 1242 3292
rect 1318 3428 1322 3432
rect 1302 3388 1306 3392
rect 1310 3358 1314 3362
rect 1294 3348 1298 3352
rect 1310 3348 1314 3352
rect 1326 3338 1330 3342
rect 1286 3308 1290 3312
rect 1326 3298 1330 3302
rect 1518 3438 1522 3442
rect 1362 3403 1366 3407
rect 1369 3403 1373 3407
rect 1342 3398 1346 3402
rect 1334 3288 1338 3292
rect 1206 3278 1210 3282
rect 1262 3278 1266 3282
rect 1406 3388 1410 3392
rect 1478 3378 1482 3382
rect 1374 3358 1378 3362
rect 1358 3348 1362 3352
rect 1374 3348 1378 3352
rect 1350 3338 1354 3342
rect 1350 3308 1354 3312
rect 1262 3268 1266 3272
rect 1310 3268 1314 3272
rect 1326 3268 1330 3272
rect 1174 3188 1178 3192
rect 982 3168 986 3172
rect 1006 3158 1010 3162
rect 918 3148 922 3152
rect 958 3148 962 3152
rect 974 3148 978 3152
rect 1006 3148 1010 3152
rect 1014 3148 1018 3152
rect 1126 3148 1130 3152
rect 1142 3148 1146 3152
rect 910 3138 914 3142
rect 934 3138 938 3142
rect 982 3138 986 3142
rect 942 3128 946 3132
rect 966 3088 970 3092
rect 910 3078 914 3082
rect 1054 3078 1058 3082
rect 1102 3108 1106 3112
rect 1086 3098 1090 3102
rect 1134 3078 1138 3082
rect 1078 3068 1082 3072
rect 1110 3068 1114 3072
rect 950 3058 954 3062
rect 1134 3058 1138 3062
rect 902 3028 906 3032
rect 1006 3048 1010 3052
rect 918 2998 922 3002
rect 958 2998 962 3002
rect 918 2968 922 2972
rect 854 2868 858 2872
rect 822 2858 826 2862
rect 838 2858 842 2862
rect 862 2858 866 2862
rect 886 2858 890 2862
rect 854 2848 858 2852
rect 838 2838 842 2842
rect 854 2808 858 2812
rect 838 2768 842 2772
rect 878 2818 882 2822
rect 822 2748 826 2752
rect 918 2958 922 2962
rect 942 2958 946 2962
rect 934 2938 938 2942
rect 902 2928 906 2932
rect 910 2918 914 2922
rect 934 2918 938 2922
rect 1086 3048 1090 3052
rect 1110 3048 1114 3052
rect 1062 3038 1066 3042
rect 1078 3038 1082 3042
rect 1030 3028 1034 3032
rect 966 2978 970 2982
rect 1006 2968 1010 2972
rect 974 2958 978 2962
rect 974 2938 978 2942
rect 982 2928 986 2932
rect 950 2908 954 2912
rect 918 2878 922 2882
rect 910 2858 914 2862
rect 894 2808 898 2812
rect 1006 2918 1010 2922
rect 990 2888 994 2892
rect 998 2888 1002 2892
rect 1134 3038 1138 3042
rect 1110 3028 1114 3032
rect 1126 3008 1130 3012
rect 1078 2998 1082 3002
rect 1222 3258 1226 3262
rect 1230 3258 1234 3262
rect 1286 3258 1290 3262
rect 1302 3258 1306 3262
rect 1262 3248 1266 3252
rect 1230 3228 1234 3232
rect 1262 3228 1266 3232
rect 1270 3228 1274 3232
rect 1302 3198 1306 3202
rect 1278 3188 1282 3192
rect 1206 3148 1210 3152
rect 1262 3148 1266 3152
rect 1198 3128 1202 3132
rect 1182 3048 1186 3052
rect 1174 3028 1178 3032
rect 1086 2928 1090 2932
rect 1054 2918 1058 2922
rect 950 2848 954 2852
rect 966 2818 970 2822
rect 918 2788 922 2792
rect 926 2768 930 2772
rect 902 2758 906 2762
rect 926 2758 930 2762
rect 942 2758 946 2762
rect 894 2748 898 2752
rect 838 2738 842 2742
rect 886 2738 890 2742
rect 830 2728 834 2732
rect 830 2708 834 2712
rect 850 2703 854 2707
rect 857 2703 861 2707
rect 878 2698 882 2702
rect 910 2738 914 2742
rect 902 2718 906 2722
rect 1006 2838 1010 2842
rect 1022 2808 1026 2812
rect 1094 2878 1098 2882
rect 1078 2858 1082 2862
rect 1046 2828 1050 2832
rect 1046 2808 1050 2812
rect 1014 2758 1018 2762
rect 1030 2758 1034 2762
rect 942 2738 946 2742
rect 950 2738 954 2742
rect 974 2738 978 2742
rect 934 2728 938 2732
rect 950 2728 954 2732
rect 990 2728 994 2732
rect 926 2698 930 2702
rect 846 2688 850 2692
rect 894 2688 898 2692
rect 918 2688 922 2692
rect 862 2678 866 2682
rect 1030 2738 1034 2742
rect 1022 2728 1026 2732
rect 1046 2728 1050 2732
rect 998 2718 1002 2722
rect 958 2708 962 2712
rect 966 2708 970 2712
rect 1046 2708 1050 2712
rect 950 2688 954 2692
rect 974 2688 978 2692
rect 998 2688 1002 2692
rect 1030 2688 1034 2692
rect 926 2678 930 2682
rect 990 2678 994 2682
rect 958 2668 962 2672
rect 830 2628 834 2632
rect 766 2618 770 2622
rect 806 2618 810 2622
rect 918 2658 922 2662
rect 950 2658 954 2662
rect 902 2648 906 2652
rect 910 2648 914 2652
rect 894 2628 898 2632
rect 846 2608 850 2612
rect 782 2588 786 2592
rect 830 2588 834 2592
rect 838 2588 842 2592
rect 710 2568 714 2572
rect 758 2568 762 2572
rect 694 2558 698 2562
rect 726 2558 730 2562
rect 758 2558 762 2562
rect 678 2548 682 2552
rect 574 2538 578 2542
rect 630 2538 634 2542
rect 558 2518 562 2522
rect 606 2528 610 2532
rect 622 2508 626 2512
rect 630 2498 634 2502
rect 638 2488 642 2492
rect 486 2478 490 2482
rect 598 2478 602 2482
rect 534 2458 538 2462
rect 494 2448 498 2452
rect 494 2428 498 2432
rect 638 2468 642 2472
rect 742 2548 746 2552
rect 734 2538 738 2542
rect 710 2518 714 2522
rect 686 2508 690 2512
rect 822 2568 826 2572
rect 798 2558 802 2562
rect 798 2548 802 2552
rect 782 2528 786 2532
rect 806 2518 810 2522
rect 830 2548 834 2552
rect 862 2598 866 2602
rect 870 2598 874 2602
rect 902 2608 906 2612
rect 886 2568 890 2572
rect 894 2558 898 2562
rect 878 2548 882 2552
rect 846 2538 850 2542
rect 822 2518 826 2522
rect 750 2508 754 2512
rect 782 2508 786 2512
rect 814 2508 818 2512
rect 670 2488 674 2492
rect 598 2438 602 2442
rect 646 2438 650 2442
rect 590 2408 594 2412
rect 550 2398 554 2402
rect 486 2378 490 2382
rect 526 2378 530 2382
rect 558 2378 562 2382
rect 542 2368 546 2372
rect 614 2378 618 2382
rect 606 2368 610 2372
rect 518 2358 522 2362
rect 622 2358 626 2362
rect 494 2348 498 2352
rect 614 2348 618 2352
rect 430 2338 434 2342
rect 446 2338 450 2342
rect 478 2338 482 2342
rect 486 2298 490 2302
rect 462 2278 466 2282
rect 414 2268 418 2272
rect 390 2258 394 2262
rect 246 2248 250 2252
rect 346 2203 350 2207
rect 353 2203 357 2207
rect 358 2158 362 2162
rect 422 2148 426 2152
rect 374 2118 378 2122
rect 238 2098 242 2102
rect 398 2108 402 2112
rect 438 2098 442 2102
rect 398 2088 402 2092
rect 478 2258 482 2262
rect 470 2208 474 2212
rect 510 2338 514 2342
rect 558 2338 562 2342
rect 526 2328 530 2332
rect 550 2298 554 2302
rect 518 2258 522 2262
rect 590 2208 594 2212
rect 654 2408 658 2412
rect 710 2478 714 2482
rect 678 2468 682 2472
rect 686 2468 690 2472
rect 670 2388 674 2392
rect 638 2378 642 2382
rect 670 2368 674 2372
rect 678 2368 682 2372
rect 702 2448 706 2452
rect 662 2348 666 2352
rect 694 2348 698 2352
rect 726 2458 730 2462
rect 742 2458 746 2462
rect 766 2458 770 2462
rect 806 2478 810 2482
rect 790 2448 794 2452
rect 782 2438 786 2442
rect 758 2378 762 2382
rect 790 2418 794 2422
rect 774 2368 778 2372
rect 718 2358 722 2362
rect 742 2348 746 2352
rect 758 2348 762 2352
rect 806 2458 810 2462
rect 894 2538 898 2542
rect 870 2508 874 2512
rect 850 2503 854 2507
rect 857 2503 861 2507
rect 830 2468 834 2472
rect 838 2458 842 2462
rect 894 2458 898 2462
rect 902 2458 906 2462
rect 870 2448 874 2452
rect 838 2428 842 2432
rect 830 2368 834 2372
rect 862 2368 866 2372
rect 830 2358 834 2362
rect 814 2348 818 2352
rect 918 2608 922 2612
rect 918 2538 922 2542
rect 918 2528 922 2532
rect 1086 2838 1090 2842
rect 1070 2818 1074 2822
rect 1062 2738 1066 2742
rect 1062 2718 1066 2722
rect 1038 2668 1042 2672
rect 1022 2658 1026 2662
rect 982 2628 986 2632
rect 1006 2628 1010 2632
rect 1014 2628 1018 2632
rect 974 2598 978 2602
rect 1046 2598 1050 2602
rect 934 2588 938 2592
rect 974 2588 978 2592
rect 974 2568 978 2572
rect 1006 2568 1010 2572
rect 950 2548 954 2552
rect 982 2548 986 2552
rect 1094 2738 1098 2742
rect 1078 2698 1082 2702
rect 1078 2678 1082 2682
rect 1086 2668 1090 2672
rect 1062 2608 1066 2612
rect 1086 2628 1090 2632
rect 1078 2598 1082 2602
rect 1078 2558 1082 2562
rect 1422 3338 1426 3342
rect 1390 3318 1394 3322
rect 1382 3288 1386 3292
rect 1334 3258 1338 3262
rect 1358 3248 1362 3252
rect 1334 3228 1338 3232
rect 1318 3138 1322 3142
rect 1246 3098 1250 3102
rect 1362 3203 1366 3207
rect 1369 3203 1373 3207
rect 1342 3198 1346 3202
rect 1262 3078 1266 3082
rect 1326 3048 1330 3052
rect 1278 2988 1282 2992
rect 1222 2968 1226 2972
rect 1262 2968 1266 2972
rect 1294 2978 1298 2982
rect 1318 2978 1322 2982
rect 1286 2968 1290 2972
rect 1206 2958 1210 2962
rect 1230 2958 1234 2962
rect 1310 2958 1314 2962
rect 1318 2958 1322 2962
rect 1350 3088 1354 3092
rect 1382 3068 1386 3072
rect 1374 3058 1378 3062
rect 1582 3398 1586 3402
rect 1614 3418 1618 3422
rect 1718 3398 1722 3402
rect 1622 3388 1626 3392
rect 1742 3378 1746 3382
rect 1590 3368 1594 3372
rect 1598 3368 1602 3372
rect 1622 3368 1626 3372
rect 1558 3348 1562 3352
rect 1598 3338 1602 3342
rect 1494 3328 1498 3332
rect 1606 3328 1610 3332
rect 1478 3318 1482 3322
rect 1590 3318 1594 3322
rect 1398 3288 1402 3292
rect 1462 3288 1466 3292
rect 1406 3278 1410 3282
rect 1510 3308 1514 3312
rect 1502 3288 1506 3292
rect 1486 3278 1490 3282
rect 1398 3248 1402 3252
rect 1406 3248 1410 3252
rect 1446 3248 1450 3252
rect 1486 3248 1490 3252
rect 1398 3208 1402 3212
rect 1454 3208 1458 3212
rect 1494 3168 1498 3172
rect 1510 3248 1514 3252
rect 1542 3238 1546 3242
rect 1550 3238 1554 3242
rect 1526 3228 1530 3232
rect 1526 3178 1530 3182
rect 1534 3168 1538 3172
rect 1414 3158 1418 3162
rect 1430 3158 1434 3162
rect 1518 3158 1522 3162
rect 1526 3158 1530 3162
rect 1422 3148 1426 3152
rect 1454 3148 1458 3152
rect 1486 3148 1490 3152
rect 1414 3138 1418 3142
rect 1462 3138 1466 3142
rect 1406 3128 1410 3132
rect 1438 3128 1442 3132
rect 1478 3128 1482 3132
rect 1454 3078 1458 3082
rect 1470 3078 1474 3082
rect 1478 3068 1482 3072
rect 1430 3058 1434 3062
rect 1454 3058 1458 3062
rect 1470 3058 1474 3062
rect 1350 3048 1354 3052
rect 1390 3048 1394 3052
rect 1398 3048 1402 3052
rect 1222 2938 1226 2942
rect 1246 2938 1250 2942
rect 1302 2938 1306 2942
rect 1190 2928 1194 2932
rect 1230 2928 1234 2932
rect 1390 3038 1394 3042
rect 1362 3003 1366 3007
rect 1369 3003 1373 3007
rect 1374 2968 1378 2972
rect 1110 2908 1114 2912
rect 1126 2908 1130 2912
rect 1142 2908 1146 2912
rect 1326 2908 1330 2912
rect 1310 2878 1314 2882
rect 1182 2868 1186 2872
rect 1270 2868 1274 2872
rect 1286 2868 1290 2872
rect 1166 2858 1170 2862
rect 1126 2788 1130 2792
rect 1270 2838 1274 2842
rect 1294 2818 1298 2822
rect 1110 2778 1114 2782
rect 1110 2758 1114 2762
rect 1214 2738 1218 2742
rect 1230 2728 1234 2732
rect 1318 2808 1322 2812
rect 1302 2798 1306 2802
rect 1334 2898 1338 2902
rect 1334 2888 1338 2892
rect 1350 2898 1354 2902
rect 1366 2898 1370 2902
rect 1358 2868 1362 2872
rect 1366 2868 1370 2872
rect 1334 2848 1338 2852
rect 1366 2848 1370 2852
rect 1334 2838 1338 2842
rect 1342 2828 1346 2832
rect 1334 2768 1338 2772
rect 1462 3038 1466 3042
rect 1422 3028 1426 3032
rect 1446 3028 1450 3032
rect 1414 3018 1418 3022
rect 1558 3208 1562 3212
rect 1510 3138 1514 3142
rect 1542 3108 1546 3112
rect 1526 3088 1530 3092
rect 1550 3088 1554 3092
rect 1534 3068 1538 3072
rect 1614 3178 1618 3182
rect 1614 3158 1618 3162
rect 1582 3138 1586 3142
rect 1574 3078 1578 3082
rect 1614 3118 1618 3122
rect 1814 3478 1818 3482
rect 1902 3508 1906 3512
rect 1882 3503 1886 3507
rect 1889 3503 1893 3507
rect 2190 3548 2194 3552
rect 1998 3538 2002 3542
rect 2014 3538 2018 3542
rect 2158 3538 2162 3542
rect 1974 3518 1978 3522
rect 1982 3508 1986 3512
rect 1950 3498 1954 3502
rect 1966 3498 1970 3502
rect 2038 3498 2042 3502
rect 1902 3468 1906 3472
rect 1862 3438 1866 3442
rect 1854 3418 1858 3422
rect 1910 3398 1914 3402
rect 2166 3528 2170 3532
rect 2190 3528 2194 3532
rect 2174 3518 2178 3522
rect 1990 3488 1994 3492
rect 2038 3488 2042 3492
rect 2094 3488 2098 3492
rect 2142 3488 2146 3492
rect 2182 3488 2186 3492
rect 2006 3458 2010 3462
rect 2046 3438 2050 3442
rect 2086 3418 2090 3422
rect 1798 3388 1802 3392
rect 2006 3388 2010 3392
rect 1982 3358 1986 3362
rect 1998 3358 2002 3362
rect 1750 3348 1754 3352
rect 1798 3348 1802 3352
rect 1678 3328 1682 3332
rect 1774 3338 1778 3342
rect 1854 3328 1858 3332
rect 1782 3318 1786 3322
rect 1694 3298 1698 3302
rect 1758 3298 1762 3302
rect 1974 3318 1978 3322
rect 1882 3303 1886 3307
rect 1889 3303 1893 3307
rect 1702 3288 1706 3292
rect 1790 3288 1794 3292
rect 1870 3288 1874 3292
rect 1630 3278 1634 3282
rect 1662 3278 1666 3282
rect 1686 3278 1690 3282
rect 1694 3278 1698 3282
rect 1638 3268 1642 3272
rect 1678 3268 1682 3272
rect 1686 3158 1690 3162
rect 1638 3148 1642 3152
rect 1654 3148 1658 3152
rect 1630 3128 1634 3132
rect 1614 3088 1618 3092
rect 1598 3078 1602 3082
rect 1630 3078 1634 3082
rect 1646 3078 1650 3082
rect 1502 3058 1506 3062
rect 1526 3058 1530 3062
rect 1542 3058 1546 3062
rect 1558 3058 1562 3062
rect 1494 3048 1498 3052
rect 1446 2978 1450 2982
rect 1486 2968 1490 2972
rect 1454 2958 1458 2962
rect 1470 2958 1474 2962
rect 1406 2938 1410 2942
rect 1422 2938 1426 2942
rect 1438 2938 1442 2942
rect 1398 2918 1402 2922
rect 1430 2868 1434 2872
rect 1398 2838 1402 2842
rect 1390 2828 1394 2832
rect 1406 2828 1410 2832
rect 1382 2808 1386 2812
rect 1362 2803 1366 2807
rect 1369 2803 1373 2807
rect 1422 2858 1426 2862
rect 1446 2858 1450 2862
rect 1462 2928 1466 2932
rect 1462 2918 1466 2922
rect 1550 3038 1554 3042
rect 1574 2998 1578 3002
rect 1590 3048 1594 3052
rect 1638 3048 1642 3052
rect 1630 3038 1634 3042
rect 1606 3028 1610 3032
rect 1630 2998 1634 3002
rect 1542 2988 1546 2992
rect 1582 2988 1586 2992
rect 1574 2968 1578 2972
rect 1622 2968 1626 2972
rect 1558 2958 1562 2962
rect 1614 2958 1618 2962
rect 1518 2938 1522 2942
rect 1470 2868 1474 2872
rect 1470 2848 1474 2852
rect 1550 2938 1554 2942
rect 1534 2918 1538 2922
rect 1494 2878 1498 2882
rect 1510 2878 1514 2882
rect 1470 2838 1474 2842
rect 1486 2838 1490 2842
rect 1454 2828 1458 2832
rect 1454 2798 1458 2802
rect 1534 2908 1538 2912
rect 1526 2828 1530 2832
rect 1486 2788 1490 2792
rect 1414 2768 1418 2772
rect 1470 2768 1474 2772
rect 1366 2758 1370 2762
rect 1478 2758 1482 2762
rect 1342 2748 1346 2752
rect 1398 2748 1402 2752
rect 1462 2748 1466 2752
rect 1406 2738 1410 2742
rect 1118 2718 1122 2722
rect 1294 2718 1298 2722
rect 1102 2668 1106 2672
rect 1102 2628 1106 2632
rect 1150 2688 1154 2692
rect 1166 2688 1170 2692
rect 1126 2678 1130 2682
rect 1142 2618 1146 2622
rect 1118 2578 1122 2582
rect 1094 2548 1098 2552
rect 1094 2538 1098 2542
rect 1134 2538 1138 2542
rect 1006 2498 1010 2502
rect 926 2488 930 2492
rect 934 2488 938 2492
rect 950 2488 954 2492
rect 998 2488 1002 2492
rect 1014 2488 1018 2492
rect 926 2468 930 2472
rect 958 2468 962 2472
rect 998 2468 1002 2472
rect 910 2448 914 2452
rect 910 2428 914 2432
rect 910 2388 914 2392
rect 934 2458 938 2462
rect 950 2458 954 2462
rect 966 2458 970 2462
rect 942 2398 946 2402
rect 918 2358 922 2362
rect 926 2358 930 2362
rect 886 2348 890 2352
rect 702 2338 706 2342
rect 718 2338 722 2342
rect 806 2338 810 2342
rect 878 2338 882 2342
rect 678 2328 682 2332
rect 686 2328 690 2332
rect 790 2328 794 2332
rect 742 2308 746 2312
rect 734 2298 738 2302
rect 758 2298 762 2302
rect 678 2268 682 2272
rect 926 2338 930 2342
rect 934 2338 938 2342
rect 902 2318 906 2322
rect 894 2308 898 2312
rect 926 2308 930 2312
rect 850 2303 854 2307
rect 857 2303 861 2307
rect 638 2258 642 2262
rect 694 2258 698 2262
rect 838 2258 842 2262
rect 862 2258 866 2262
rect 894 2258 898 2262
rect 638 2238 642 2242
rect 630 2188 634 2192
rect 566 2178 570 2182
rect 598 2178 602 2182
rect 630 2178 634 2182
rect 526 2168 530 2172
rect 550 2168 554 2172
rect 542 2158 546 2162
rect 462 2148 466 2152
rect 518 2148 522 2152
rect 454 2138 458 2142
rect 222 2078 226 2082
rect 262 2078 266 2082
rect 414 2078 418 2082
rect 446 2078 450 2082
rect 270 2068 274 2072
rect 358 2068 362 2072
rect 62 2058 66 2062
rect 86 2058 90 2062
rect 326 2058 330 2062
rect 86 2048 90 2052
rect 94 2028 98 2032
rect 134 2018 138 2022
rect 38 2008 42 2012
rect 14 1988 18 1992
rect 30 1978 34 1982
rect 22 1958 26 1962
rect 70 1958 74 1962
rect 318 2048 322 2052
rect 294 2018 298 2022
rect 270 2008 274 2012
rect 286 1968 290 1972
rect 38 1948 42 1952
rect 54 1948 58 1952
rect 70 1948 74 1952
rect 254 1948 258 1952
rect 346 2003 350 2007
rect 353 2003 357 2007
rect 318 1998 322 2002
rect 270 1938 274 1942
rect 310 1938 314 1942
rect 358 1968 362 1972
rect 374 1968 378 1972
rect 390 1968 394 1972
rect 190 1928 194 1932
rect 318 1928 322 1932
rect 174 1918 178 1922
rect 262 1918 266 1922
rect 30 1908 34 1912
rect 94 1898 98 1902
rect 222 1898 226 1902
rect 150 1878 154 1882
rect 134 1868 138 1872
rect 206 1858 210 1862
rect 246 1858 250 1862
rect 230 1788 234 1792
rect 6 1748 10 1752
rect 190 1748 194 1752
rect 206 1748 210 1752
rect 134 1728 138 1732
rect 118 1718 122 1722
rect 94 1668 98 1672
rect 302 1898 306 1902
rect 334 1908 338 1912
rect 366 1878 370 1882
rect 374 1868 378 1872
rect 366 1858 370 1862
rect 302 1848 306 1852
rect 346 1803 350 1807
rect 353 1803 357 1807
rect 326 1768 330 1772
rect 366 1768 370 1772
rect 358 1758 362 1762
rect 302 1748 306 1752
rect 326 1748 330 1752
rect 342 1748 346 1752
rect 310 1738 314 1742
rect 334 1738 338 1742
rect 286 1728 290 1732
rect 358 1728 362 1732
rect 270 1708 274 1712
rect 246 1678 250 1682
rect 214 1668 218 1672
rect 110 1658 114 1662
rect 166 1658 170 1662
rect 206 1658 210 1662
rect 14 1588 18 1592
rect 30 1578 34 1582
rect 190 1578 194 1582
rect 126 1538 130 1542
rect 158 1538 162 1542
rect 62 1508 66 1512
rect 86 1508 90 1512
rect 46 1498 50 1502
rect 366 1668 370 1672
rect 302 1658 306 1662
rect 334 1658 338 1662
rect 294 1558 298 1562
rect 318 1558 322 1562
rect 326 1538 330 1542
rect 294 1528 298 1532
rect 262 1508 266 1512
rect 302 1498 306 1502
rect 158 1488 162 1492
rect 206 1488 210 1492
rect 262 1488 266 1492
rect 14 1448 18 1452
rect 70 1408 74 1412
rect 46 1388 50 1392
rect 30 1338 34 1342
rect 302 1468 306 1472
rect 206 1448 210 1452
rect 246 1448 250 1452
rect 174 1418 178 1422
rect 174 1328 178 1332
rect 118 1318 122 1322
rect 38 1278 42 1282
rect 110 1268 114 1272
rect 158 1268 162 1272
rect 166 1268 170 1272
rect 6 1048 10 1052
rect 30 1078 34 1082
rect 30 1058 34 1062
rect 254 1408 258 1412
rect 270 1368 274 1372
rect 294 1368 298 1372
rect 254 1348 258 1352
rect 278 1348 282 1352
rect 222 1328 226 1332
rect 206 1268 210 1272
rect 222 1248 226 1252
rect 182 1238 186 1242
rect 206 1238 210 1242
rect 86 1198 90 1202
rect 118 1198 122 1202
rect 270 1288 274 1292
rect 254 1218 258 1222
rect 214 1188 218 1192
rect 254 1188 258 1192
rect 310 1358 314 1362
rect 302 1248 306 1252
rect 278 1168 282 1172
rect 182 1148 186 1152
rect 286 1148 290 1152
rect 70 1128 74 1132
rect 134 1088 138 1092
rect 254 1138 258 1142
rect 222 1108 226 1112
rect 238 1088 242 1092
rect 190 1078 194 1082
rect 230 1078 234 1082
rect 350 1628 354 1632
rect 346 1603 350 1607
rect 353 1603 357 1607
rect 342 1548 346 1552
rect 486 2058 490 2062
rect 502 2128 506 2132
rect 510 2128 514 2132
rect 502 2088 506 2092
rect 502 2078 506 2082
rect 526 2068 530 2072
rect 494 2038 498 2042
rect 526 2008 530 2012
rect 510 1988 514 1992
rect 518 1958 522 1962
rect 462 1918 466 1922
rect 446 1908 450 1912
rect 462 1908 466 1912
rect 406 1858 410 1862
rect 406 1818 410 1822
rect 438 1778 442 1782
rect 470 1878 474 1882
rect 494 1898 498 1902
rect 566 2158 570 2162
rect 590 2158 594 2162
rect 622 2158 626 2162
rect 566 2118 570 2122
rect 630 2148 634 2152
rect 590 2128 594 2132
rect 662 2228 666 2232
rect 662 2178 666 2182
rect 646 2128 650 2132
rect 654 2078 658 2082
rect 630 2058 634 2062
rect 598 2048 602 2052
rect 590 2038 594 2042
rect 590 2028 594 2032
rect 598 2028 602 2032
rect 582 2018 586 2022
rect 574 1998 578 2002
rect 574 1978 578 1982
rect 558 1948 562 1952
rect 598 1998 602 2002
rect 550 1938 554 1942
rect 566 1938 570 1942
rect 582 1938 586 1942
rect 582 1908 586 1912
rect 590 1898 594 1902
rect 590 1888 594 1892
rect 558 1878 562 1882
rect 566 1878 570 1882
rect 654 2008 658 2012
rect 638 1968 642 1972
rect 614 1958 618 1962
rect 638 1958 642 1962
rect 606 1878 610 1882
rect 462 1858 466 1862
rect 550 1858 554 1862
rect 630 1948 634 1952
rect 646 1948 650 1952
rect 622 1918 626 1922
rect 686 2148 690 2152
rect 670 2098 674 2102
rect 678 2038 682 2042
rect 670 2008 674 2012
rect 662 1968 666 1972
rect 910 2248 914 2252
rect 758 2208 762 2212
rect 822 2188 826 2192
rect 710 2168 714 2172
rect 774 2168 778 2172
rect 742 2158 746 2162
rect 758 2158 762 2162
rect 806 2158 810 2162
rect 862 2198 866 2202
rect 838 2178 842 2182
rect 718 2148 722 2152
rect 798 2148 802 2152
rect 886 2148 890 2152
rect 758 2138 762 2142
rect 822 2138 826 2142
rect 870 2138 874 2142
rect 814 2128 818 2132
rect 758 2108 762 2112
rect 814 2108 818 2112
rect 806 2068 810 2072
rect 742 2058 746 2062
rect 798 2048 802 2052
rect 694 2018 698 2022
rect 742 2018 746 2022
rect 694 2008 698 2012
rect 710 2008 714 2012
rect 702 1988 706 1992
rect 694 1968 698 1972
rect 686 1958 690 1962
rect 670 1948 674 1952
rect 718 1948 722 1952
rect 678 1938 682 1942
rect 694 1938 698 1942
rect 702 1928 706 1932
rect 726 1928 730 1932
rect 678 1878 682 1882
rect 774 1998 778 2002
rect 798 1998 802 2002
rect 850 2103 854 2107
rect 857 2103 861 2107
rect 950 2368 954 2372
rect 1014 2478 1018 2482
rect 1038 2478 1042 2482
rect 1030 2458 1034 2462
rect 1062 2528 1066 2532
rect 1126 2528 1130 2532
rect 1078 2518 1082 2522
rect 1126 2518 1130 2522
rect 1062 2508 1066 2512
rect 1094 2508 1098 2512
rect 1094 2488 1098 2492
rect 1118 2488 1122 2492
rect 1086 2468 1090 2472
rect 1054 2438 1058 2442
rect 1014 2398 1018 2402
rect 1030 2378 1034 2382
rect 1078 2358 1082 2362
rect 998 2348 1002 2352
rect 1070 2348 1074 2352
rect 974 2318 978 2322
rect 1022 2298 1026 2302
rect 1014 2288 1018 2292
rect 950 2268 954 2272
rect 958 2268 962 2272
rect 982 2268 986 2272
rect 1006 2258 1010 2262
rect 1046 2318 1050 2322
rect 1070 2278 1074 2282
rect 1118 2448 1122 2452
rect 1150 2568 1154 2572
rect 1222 2668 1226 2672
rect 1238 2658 1242 2662
rect 1294 2658 1298 2662
rect 1222 2648 1226 2652
rect 1310 2678 1314 2682
rect 1182 2638 1186 2642
rect 1302 2648 1306 2652
rect 1294 2638 1298 2642
rect 1294 2608 1298 2612
rect 1246 2598 1250 2602
rect 1206 2568 1210 2572
rect 1270 2558 1274 2562
rect 1230 2548 1234 2552
rect 1182 2538 1186 2542
rect 1198 2538 1202 2542
rect 1214 2528 1218 2532
rect 1246 2538 1250 2542
rect 1262 2538 1266 2542
rect 1230 2528 1234 2532
rect 1158 2518 1162 2522
rect 1198 2518 1202 2522
rect 1238 2508 1242 2512
rect 1214 2488 1218 2492
rect 1270 2528 1274 2532
rect 1286 2508 1290 2512
rect 1166 2478 1170 2482
rect 1206 2478 1210 2482
rect 1246 2478 1250 2482
rect 1158 2468 1162 2472
rect 1150 2458 1154 2462
rect 1110 2438 1114 2442
rect 1126 2438 1130 2442
rect 1142 2418 1146 2422
rect 1134 2388 1138 2392
rect 1206 2458 1210 2462
rect 1206 2448 1210 2452
rect 1230 2438 1234 2442
rect 1182 2428 1186 2432
rect 1222 2428 1226 2432
rect 1174 2408 1178 2412
rect 1222 2408 1226 2412
rect 1206 2348 1210 2352
rect 1094 2298 1098 2302
rect 1062 2258 1066 2262
rect 1086 2258 1090 2262
rect 1078 2248 1082 2252
rect 1110 2288 1114 2292
rect 1102 2278 1106 2282
rect 1118 2278 1122 2282
rect 1190 2318 1194 2322
rect 1270 2438 1274 2442
rect 1310 2458 1314 2462
rect 1286 2418 1290 2422
rect 1278 2408 1282 2412
rect 1254 2398 1258 2402
rect 1294 2398 1298 2402
rect 1270 2358 1274 2362
rect 1334 2658 1338 2662
rect 1438 2738 1442 2742
rect 1422 2708 1426 2712
rect 1350 2698 1354 2702
rect 1390 2678 1394 2682
rect 1406 2668 1410 2672
rect 1446 2668 1450 2672
rect 1362 2603 1366 2607
rect 1369 2603 1373 2607
rect 1342 2568 1346 2572
rect 1382 2558 1386 2562
rect 1342 2518 1346 2522
rect 1318 2438 1322 2442
rect 1362 2403 1366 2407
rect 1369 2403 1373 2407
rect 1326 2398 1330 2402
rect 1310 2358 1314 2362
rect 1382 2358 1386 2362
rect 1366 2348 1370 2352
rect 1246 2338 1250 2342
rect 1174 2288 1178 2292
rect 1222 2288 1226 2292
rect 1110 2258 1114 2262
rect 1150 2258 1154 2262
rect 1030 2238 1034 2242
rect 990 2218 994 2222
rect 990 2198 994 2202
rect 1134 2238 1138 2242
rect 1158 2238 1162 2242
rect 1134 2228 1138 2232
rect 1102 2168 1106 2172
rect 1126 2168 1130 2172
rect 958 2148 962 2152
rect 1014 2148 1018 2152
rect 1110 2158 1114 2162
rect 1134 2158 1138 2162
rect 1038 2138 1042 2142
rect 1046 2138 1050 2142
rect 1126 2138 1130 2142
rect 1150 2138 1154 2142
rect 958 2118 962 2122
rect 942 2108 946 2112
rect 886 2078 890 2082
rect 918 2078 922 2082
rect 886 2058 890 2062
rect 742 1928 746 1932
rect 814 1918 818 1922
rect 774 1908 778 1912
rect 806 1908 810 1912
rect 638 1858 642 1862
rect 454 1848 458 1852
rect 494 1848 498 1852
rect 598 1848 602 1852
rect 462 1838 466 1842
rect 486 1828 490 1832
rect 486 1818 490 1822
rect 470 1798 474 1802
rect 446 1758 450 1762
rect 462 1748 466 1752
rect 478 1748 482 1752
rect 526 1808 530 1812
rect 550 1808 554 1812
rect 518 1778 522 1782
rect 502 1768 506 1772
rect 526 1768 530 1772
rect 494 1748 498 1752
rect 582 1838 586 1842
rect 566 1828 570 1832
rect 614 1818 618 1822
rect 582 1808 586 1812
rect 574 1778 578 1782
rect 566 1768 570 1772
rect 542 1748 546 1752
rect 558 1748 562 1752
rect 422 1738 426 1742
rect 406 1698 410 1702
rect 382 1568 386 1572
rect 430 1728 434 1732
rect 534 1738 538 1742
rect 486 1718 490 1722
rect 486 1708 490 1712
rect 446 1698 450 1702
rect 494 1698 498 1702
rect 526 1728 530 1732
rect 574 1718 578 1722
rect 438 1688 442 1692
rect 486 1688 490 1692
rect 742 1858 746 1862
rect 654 1848 658 1852
rect 678 1848 682 1852
rect 646 1828 650 1832
rect 630 1798 634 1802
rect 646 1768 650 1772
rect 718 1848 722 1852
rect 702 1828 706 1832
rect 686 1788 690 1792
rect 686 1768 690 1772
rect 694 1768 698 1772
rect 590 1758 594 1762
rect 662 1758 666 1762
rect 638 1748 642 1752
rect 654 1738 658 1742
rect 678 1748 682 1752
rect 670 1738 674 1742
rect 662 1728 666 1732
rect 678 1728 682 1732
rect 622 1718 626 1722
rect 630 1718 634 1722
rect 598 1698 602 1702
rect 606 1678 610 1682
rect 622 1668 626 1672
rect 438 1658 442 1662
rect 542 1658 546 1662
rect 510 1618 514 1622
rect 454 1598 458 1602
rect 470 1588 474 1592
rect 438 1558 442 1562
rect 494 1558 498 1562
rect 414 1548 418 1552
rect 462 1548 466 1552
rect 398 1538 402 1542
rect 438 1538 442 1542
rect 454 1538 458 1542
rect 382 1508 386 1512
rect 446 1528 450 1532
rect 406 1498 410 1502
rect 382 1488 386 1492
rect 390 1488 394 1492
rect 398 1478 402 1482
rect 438 1498 442 1502
rect 422 1478 426 1482
rect 414 1468 418 1472
rect 430 1468 434 1472
rect 406 1448 410 1452
rect 430 1438 434 1442
rect 414 1428 418 1432
rect 346 1403 350 1407
rect 353 1403 357 1407
rect 494 1518 498 1522
rect 518 1538 522 1542
rect 510 1508 514 1512
rect 574 1648 578 1652
rect 598 1658 602 1662
rect 590 1628 594 1632
rect 574 1618 578 1622
rect 638 1688 642 1692
rect 694 1718 698 1722
rect 710 1698 714 1702
rect 646 1668 650 1672
rect 686 1668 690 1672
rect 662 1658 666 1662
rect 654 1648 658 1652
rect 710 1648 714 1652
rect 606 1628 610 1632
rect 598 1608 602 1612
rect 550 1588 554 1592
rect 590 1578 594 1582
rect 558 1568 562 1572
rect 574 1568 578 1572
rect 614 1598 618 1602
rect 582 1548 586 1552
rect 646 1568 650 1572
rect 686 1638 690 1642
rect 766 1848 770 1852
rect 734 1818 738 1822
rect 758 1758 762 1762
rect 750 1748 754 1752
rect 766 1738 770 1742
rect 758 1728 762 1732
rect 750 1718 754 1722
rect 758 1718 762 1722
rect 734 1708 738 1712
rect 726 1658 730 1662
rect 718 1608 722 1612
rect 670 1578 674 1582
rect 694 1578 698 1582
rect 678 1568 682 1572
rect 694 1568 698 1572
rect 718 1568 722 1572
rect 574 1538 578 1542
rect 590 1538 594 1542
rect 606 1538 610 1542
rect 638 1528 642 1532
rect 622 1518 626 1522
rect 462 1488 466 1492
rect 526 1488 530 1492
rect 478 1478 482 1482
rect 526 1478 530 1482
rect 534 1478 538 1482
rect 486 1468 490 1472
rect 454 1438 458 1442
rect 446 1428 450 1432
rect 438 1408 442 1412
rect 382 1398 386 1402
rect 374 1388 378 1392
rect 334 1378 338 1382
rect 334 1328 338 1332
rect 398 1318 402 1322
rect 446 1298 450 1302
rect 398 1278 402 1282
rect 342 1268 346 1272
rect 382 1268 386 1272
rect 374 1218 378 1222
rect 454 1218 458 1222
rect 346 1203 350 1207
rect 353 1203 357 1207
rect 286 1138 290 1142
rect 342 1138 346 1142
rect 278 1128 282 1132
rect 262 1108 266 1112
rect 278 1098 282 1102
rect 54 1058 58 1062
rect 230 1058 234 1062
rect 246 1058 250 1062
rect 262 1018 266 1022
rect 118 978 122 982
rect 14 918 18 922
rect 238 988 242 992
rect 238 968 242 972
rect 310 1118 314 1122
rect 326 1108 330 1112
rect 318 1098 322 1102
rect 310 1088 314 1092
rect 294 1058 298 1062
rect 342 1118 346 1122
rect 334 1088 338 1092
rect 318 1058 322 1062
rect 302 1048 306 1052
rect 310 1048 314 1052
rect 318 1048 322 1052
rect 346 1003 350 1007
rect 353 1003 357 1007
rect 470 1448 474 1452
rect 486 1448 490 1452
rect 518 1408 522 1412
rect 494 1368 498 1372
rect 502 1368 506 1372
rect 670 1488 674 1492
rect 614 1478 618 1482
rect 630 1468 634 1472
rect 574 1438 578 1442
rect 550 1398 554 1402
rect 598 1398 602 1402
rect 662 1388 666 1392
rect 646 1378 650 1382
rect 558 1368 562 1372
rect 582 1368 586 1372
rect 542 1358 546 1362
rect 510 1348 514 1352
rect 526 1338 530 1342
rect 470 1288 474 1292
rect 502 1278 506 1282
rect 478 1268 482 1272
rect 502 1258 506 1262
rect 598 1348 602 1352
rect 542 1338 546 1342
rect 558 1328 562 1332
rect 542 1318 546 1322
rect 534 1308 538 1312
rect 534 1298 538 1302
rect 590 1338 594 1342
rect 582 1308 586 1312
rect 518 1268 522 1272
rect 566 1268 570 1272
rect 430 1168 434 1172
rect 478 1168 482 1172
rect 502 1168 506 1172
rect 526 1168 530 1172
rect 542 1168 546 1172
rect 510 1158 514 1162
rect 430 1148 434 1152
rect 438 1148 442 1152
rect 454 1148 458 1152
rect 478 1148 482 1152
rect 494 1148 498 1152
rect 542 1148 546 1152
rect 446 1138 450 1142
rect 550 1138 554 1142
rect 454 1118 458 1122
rect 470 1118 474 1122
rect 422 1108 426 1112
rect 462 1098 466 1102
rect 454 1088 458 1092
rect 438 1068 442 1072
rect 454 1038 458 1042
rect 438 1028 442 1032
rect 422 998 426 1002
rect 302 978 306 982
rect 390 978 394 982
rect 326 968 330 972
rect 294 958 298 962
rect 318 948 322 952
rect 334 948 338 952
rect 270 938 274 942
rect 310 938 314 942
rect 102 928 106 932
rect 46 918 50 922
rect 118 898 122 902
rect 198 898 202 902
rect 86 888 90 892
rect 238 908 242 912
rect 214 878 218 882
rect 70 858 74 862
rect 182 838 186 842
rect 174 818 178 822
rect 182 778 186 782
rect 230 848 234 852
rect 262 838 266 842
rect 254 818 258 822
rect 206 778 210 782
rect 54 768 58 772
rect 126 768 130 772
rect 158 768 162 772
rect 198 768 202 772
rect 78 748 82 752
rect 102 738 106 742
rect 78 728 82 732
rect 134 748 138 752
rect 166 748 170 752
rect 150 738 154 742
rect 150 728 154 732
rect 70 698 74 702
rect 86 698 90 702
rect 86 688 90 692
rect 174 678 178 682
rect 214 748 218 752
rect 278 868 282 872
rect 310 888 314 892
rect 334 888 338 892
rect 302 868 306 872
rect 390 938 394 942
rect 382 878 386 882
rect 326 858 330 862
rect 342 858 346 862
rect 302 778 306 782
rect 310 768 314 772
rect 270 748 274 752
rect 286 748 290 752
rect 294 748 298 752
rect 302 748 306 752
rect 230 738 234 742
rect 246 728 250 732
rect 214 718 218 722
rect 230 708 234 712
rect 246 718 250 722
rect 262 718 266 722
rect 190 678 194 682
rect 198 678 202 682
rect 206 668 210 672
rect 206 658 210 662
rect 206 578 210 582
rect 14 528 18 532
rect 214 568 218 572
rect 182 548 186 552
rect 70 518 74 522
rect 86 518 90 522
rect 238 688 242 692
rect 254 698 258 702
rect 238 668 242 672
rect 278 728 282 732
rect 278 668 282 672
rect 246 568 250 572
rect 230 538 234 542
rect 222 518 226 522
rect 214 508 218 512
rect 206 498 210 502
rect 70 488 74 492
rect 174 488 178 492
rect 222 488 226 492
rect 230 488 234 492
rect 254 508 258 512
rect 246 478 250 482
rect 86 468 90 472
rect 174 468 178 472
rect 278 588 282 592
rect 286 558 290 562
rect 318 728 322 732
rect 310 688 314 692
rect 430 928 434 932
rect 406 918 410 922
rect 510 1048 514 1052
rect 486 1018 490 1022
rect 470 958 474 962
rect 494 958 498 962
rect 478 948 482 952
rect 558 1118 562 1122
rect 590 1298 594 1302
rect 582 1288 586 1292
rect 582 1238 586 1242
rect 582 1198 586 1202
rect 622 1338 626 1342
rect 686 1558 690 1562
rect 678 1368 682 1372
rect 702 1548 706 1552
rect 710 1528 714 1532
rect 742 1678 746 1682
rect 742 1668 746 1672
rect 766 1688 770 1692
rect 902 2038 906 2042
rect 894 2028 898 2032
rect 878 1998 882 2002
rect 862 1918 866 1922
rect 850 1903 854 1907
rect 857 1903 861 1907
rect 822 1878 826 1882
rect 838 1878 842 1882
rect 782 1868 786 1872
rect 790 1858 794 1862
rect 790 1848 794 1852
rect 854 1848 858 1852
rect 814 1838 818 1842
rect 806 1828 810 1832
rect 798 1788 802 1792
rect 822 1798 826 1802
rect 910 1958 914 1962
rect 950 2088 954 2092
rect 1134 2088 1138 2092
rect 1174 2278 1178 2282
rect 1198 2248 1202 2252
rect 1206 2238 1210 2242
rect 1310 2338 1314 2342
rect 1326 2338 1330 2342
rect 1334 2338 1338 2342
rect 1270 2328 1274 2332
rect 1286 2328 1290 2332
rect 1342 2328 1346 2332
rect 1278 2308 1282 2312
rect 1318 2278 1322 2282
rect 1246 2268 1250 2272
rect 1382 2338 1386 2342
rect 1374 2318 1378 2322
rect 1374 2308 1378 2312
rect 1382 2308 1386 2312
rect 1406 2488 1410 2492
rect 1438 2468 1442 2472
rect 1406 2458 1410 2462
rect 1430 2458 1434 2462
rect 1422 2428 1426 2432
rect 1486 2738 1490 2742
rect 1494 2688 1498 2692
rect 1478 2598 1482 2602
rect 1518 2808 1522 2812
rect 1510 2728 1514 2732
rect 1526 2718 1530 2722
rect 1694 3138 1698 3142
rect 1694 3098 1698 3102
rect 1678 3088 1682 3092
rect 1662 3078 1666 3082
rect 1710 3208 1714 3212
rect 1766 3208 1770 3212
rect 1726 3188 1730 3192
rect 1710 3158 1714 3162
rect 1734 3118 1738 3122
rect 1806 3198 1810 3202
rect 2086 3388 2090 3392
rect 2014 3308 2018 3312
rect 1902 3268 1906 3272
rect 1870 3248 1874 3252
rect 1886 3248 1890 3252
rect 1886 3198 1890 3202
rect 1830 3188 1834 3192
rect 1846 3188 1850 3192
rect 1790 3168 1794 3172
rect 1798 3168 1802 3172
rect 1814 3158 1818 3162
rect 1782 3138 1786 3142
rect 1782 3128 1786 3132
rect 1798 3128 1802 3132
rect 1750 3108 1754 3112
rect 1758 3108 1762 3112
rect 1734 3078 1738 3082
rect 1670 3068 1674 3072
rect 1710 3068 1714 3072
rect 1686 3058 1690 3062
rect 1742 3058 1746 3062
rect 1662 2988 1666 2992
rect 1590 2938 1594 2942
rect 1606 2938 1610 2942
rect 1566 2918 1570 2922
rect 1638 2898 1642 2902
rect 1670 2978 1674 2982
rect 1718 3018 1722 3022
rect 1678 2958 1682 2962
rect 1670 2928 1674 2932
rect 1622 2858 1626 2862
rect 1614 2758 1618 2762
rect 1550 2738 1554 2742
rect 1534 2688 1538 2692
rect 1694 2948 1698 2952
rect 1702 2898 1706 2902
rect 1718 2958 1722 2962
rect 1726 2948 1730 2952
rect 1694 2868 1698 2872
rect 1726 2868 1730 2872
rect 1822 3098 1826 3102
rect 1870 3158 1874 3162
rect 2150 3448 2154 3452
rect 2166 3448 2170 3452
rect 2198 3468 2202 3472
rect 2366 3558 2370 3562
rect 2406 3558 2410 3562
rect 2454 3568 2458 3572
rect 2478 3568 2482 3572
rect 2446 3558 2450 3562
rect 2470 3558 2474 3562
rect 2766 3578 2770 3582
rect 2750 3558 2754 3562
rect 2422 3548 2426 3552
rect 2510 3548 2514 3552
rect 2278 3538 2282 3542
rect 2358 3538 2362 3542
rect 2382 3538 2386 3542
rect 2262 3528 2266 3532
rect 2230 3508 2234 3512
rect 2246 3508 2250 3512
rect 2254 3488 2258 3492
rect 2430 3518 2434 3522
rect 2278 3508 2282 3512
rect 2270 3488 2274 3492
rect 2470 3538 2474 3542
rect 2630 3538 2634 3542
rect 2702 3538 2706 3542
rect 2494 3528 2498 3532
rect 2574 3528 2578 3532
rect 2438 3508 2442 3512
rect 2462 3508 2466 3512
rect 2526 3508 2530 3512
rect 2438 3498 2442 3502
rect 2670 3508 2674 3512
rect 2590 3498 2594 3502
rect 2566 3488 2570 3492
rect 2238 3468 2242 3472
rect 2302 3468 2306 3472
rect 2190 3458 2194 3462
rect 2222 3458 2226 3462
rect 2254 3458 2258 3462
rect 2270 3458 2274 3462
rect 2190 3448 2194 3452
rect 2214 3448 2218 3452
rect 2182 3408 2186 3412
rect 2302 3418 2306 3422
rect 2294 3388 2298 3392
rect 2174 3348 2178 3352
rect 2110 3328 2114 3332
rect 2094 3278 2098 3282
rect 2126 3268 2130 3272
rect 1926 3198 1930 3202
rect 2022 3198 2026 3202
rect 2038 3198 2042 3202
rect 2102 3198 2106 3202
rect 1934 3168 1938 3172
rect 1966 3168 1970 3172
rect 1998 3168 2002 3172
rect 2110 3168 2114 3172
rect 1902 3158 1906 3162
rect 1838 3148 1842 3152
rect 1958 3148 1962 3152
rect 2062 3158 2066 3162
rect 2086 3158 2090 3162
rect 1974 3148 1978 3152
rect 1990 3148 1994 3152
rect 1894 3138 1898 3142
rect 1926 3138 1930 3142
rect 1838 3128 1842 3132
rect 1882 3103 1886 3107
rect 1889 3103 1893 3107
rect 1870 3088 1874 3092
rect 1790 3048 1794 3052
rect 1766 3038 1770 3042
rect 1790 2998 1794 3002
rect 1886 3038 1890 3042
rect 1782 2988 1786 2992
rect 1830 2988 1834 2992
rect 1838 2928 1842 2932
rect 1742 2908 1746 2912
rect 1882 2903 1886 2907
rect 1889 2903 1893 2907
rect 1822 2898 1826 2902
rect 1854 2898 1858 2902
rect 1750 2878 1754 2882
rect 1678 2798 1682 2802
rect 1766 2858 1770 2862
rect 1742 2828 1746 2832
rect 1758 2808 1762 2812
rect 1854 2848 1858 2852
rect 1798 2818 1802 2822
rect 1758 2798 1762 2802
rect 1766 2798 1770 2802
rect 1734 2788 1738 2792
rect 1710 2778 1714 2782
rect 1726 2768 1730 2772
rect 1726 2758 1730 2762
rect 1678 2748 1682 2752
rect 1694 2748 1698 2752
rect 1750 2748 1754 2752
rect 1566 2688 1570 2692
rect 1574 2678 1578 2682
rect 1558 2668 1562 2672
rect 1582 2668 1586 2672
rect 1510 2658 1514 2662
rect 1558 2658 1562 2662
rect 1550 2618 1554 2622
rect 1542 2598 1546 2602
rect 1502 2578 1506 2582
rect 1518 2578 1522 2582
rect 1702 2738 1706 2742
rect 1694 2728 1698 2732
rect 1686 2718 1690 2722
rect 1782 2768 1786 2772
rect 1846 2798 1850 2802
rect 1854 2798 1858 2802
rect 1822 2788 1826 2792
rect 1838 2788 1842 2792
rect 1726 2708 1730 2712
rect 1630 2698 1634 2702
rect 1614 2668 1618 2672
rect 1598 2628 1602 2632
rect 1582 2608 1586 2612
rect 1646 2688 1650 2692
rect 1670 2688 1674 2692
rect 1726 2688 1730 2692
rect 1758 2688 1762 2692
rect 1654 2668 1658 2672
rect 1638 2658 1642 2662
rect 1678 2678 1682 2682
rect 1694 2678 1698 2682
rect 1686 2668 1690 2672
rect 1718 2668 1722 2672
rect 1702 2648 1706 2652
rect 1662 2628 1666 2632
rect 1782 2708 1786 2712
rect 1790 2698 1794 2702
rect 1806 2728 1810 2732
rect 1814 2728 1818 2732
rect 1854 2758 1858 2762
rect 1846 2738 1850 2742
rect 1862 2708 1866 2712
rect 1862 2698 1866 2702
rect 1742 2668 1746 2672
rect 1798 2668 1802 2672
rect 1734 2648 1738 2652
rect 1734 2628 1738 2632
rect 1726 2608 1730 2612
rect 1614 2598 1618 2602
rect 1598 2588 1602 2592
rect 1758 2658 1762 2662
rect 1750 2578 1754 2582
rect 1518 2558 1522 2562
rect 1502 2538 1506 2542
rect 1510 2538 1514 2542
rect 1526 2488 1530 2492
rect 1518 2478 1522 2482
rect 1502 2468 1506 2472
rect 1550 2538 1554 2542
rect 1542 2528 1546 2532
rect 1782 2648 1786 2652
rect 1766 2558 1770 2562
rect 1574 2548 1578 2552
rect 1774 2548 1778 2552
rect 1766 2538 1770 2542
rect 1590 2498 1594 2502
rect 1542 2448 1546 2452
rect 1534 2438 1538 2442
rect 1494 2418 1498 2422
rect 1558 2438 1562 2442
rect 1470 2408 1474 2412
rect 1550 2408 1554 2412
rect 1582 2418 1586 2422
rect 1542 2378 1546 2382
rect 1574 2378 1578 2382
rect 1414 2348 1418 2352
rect 1478 2328 1482 2332
rect 1518 2328 1522 2332
rect 1390 2298 1394 2302
rect 1462 2298 1466 2302
rect 1302 2258 1306 2262
rect 1366 2258 1370 2262
rect 1222 2188 1226 2192
rect 1230 2188 1234 2192
rect 1182 2178 1186 2182
rect 1214 2178 1218 2182
rect 1174 2138 1178 2142
rect 1190 2138 1194 2142
rect 1206 2138 1210 2142
rect 1198 2108 1202 2112
rect 1190 2088 1194 2092
rect 1030 2078 1034 2082
rect 1126 2078 1130 2082
rect 1142 2078 1146 2082
rect 1046 2068 1050 2072
rect 982 2048 986 2052
rect 934 1968 938 1972
rect 902 1918 906 1922
rect 950 2028 954 2032
rect 950 1998 954 2002
rect 1014 2008 1018 2012
rect 1030 1998 1034 2002
rect 1070 1998 1074 2002
rect 1246 2238 1250 2242
rect 1238 2108 1242 2112
rect 1230 2098 1234 2102
rect 1150 2058 1154 2062
rect 1214 2058 1218 2062
rect 1142 2048 1146 2052
rect 1078 1988 1082 1992
rect 1102 1978 1106 1982
rect 1134 1978 1138 1982
rect 958 1968 962 1972
rect 1070 1968 1074 1972
rect 1126 1968 1130 1972
rect 990 1958 994 1962
rect 1054 1958 1058 1962
rect 982 1948 986 1952
rect 950 1918 954 1922
rect 942 1908 946 1912
rect 902 1898 906 1902
rect 934 1878 938 1882
rect 894 1858 898 1862
rect 926 1868 930 1872
rect 870 1848 874 1852
rect 918 1848 922 1852
rect 902 1838 906 1842
rect 910 1828 914 1832
rect 958 1898 962 1902
rect 958 1868 962 1872
rect 958 1848 962 1852
rect 942 1808 946 1812
rect 902 1798 906 1802
rect 1014 1938 1018 1942
rect 1014 1928 1018 1932
rect 1006 1898 1010 1902
rect 998 1868 1002 1872
rect 982 1858 986 1862
rect 990 1838 994 1842
rect 998 1828 1002 1832
rect 974 1788 978 1792
rect 798 1768 802 1772
rect 854 1768 858 1772
rect 790 1758 794 1762
rect 782 1738 786 1742
rect 790 1728 794 1732
rect 774 1678 778 1682
rect 790 1678 794 1682
rect 766 1658 770 1662
rect 734 1648 738 1652
rect 750 1648 754 1652
rect 758 1608 762 1612
rect 750 1578 754 1582
rect 734 1548 738 1552
rect 822 1758 826 1762
rect 846 1758 850 1762
rect 814 1708 818 1712
rect 830 1748 834 1752
rect 830 1718 834 1722
rect 830 1708 834 1712
rect 806 1658 810 1662
rect 850 1703 854 1707
rect 857 1703 861 1707
rect 918 1778 922 1782
rect 990 1778 994 1782
rect 982 1768 986 1772
rect 998 1758 1002 1762
rect 878 1748 882 1752
rect 982 1748 986 1752
rect 918 1738 922 1742
rect 878 1718 882 1722
rect 870 1698 874 1702
rect 838 1668 842 1672
rect 838 1628 842 1632
rect 822 1578 826 1582
rect 870 1568 874 1572
rect 822 1548 826 1552
rect 742 1528 746 1532
rect 750 1518 754 1522
rect 718 1508 722 1512
rect 726 1508 730 1512
rect 726 1498 730 1502
rect 742 1448 746 1452
rect 726 1418 730 1422
rect 726 1378 730 1382
rect 710 1368 714 1372
rect 766 1508 770 1512
rect 798 1528 802 1532
rect 838 1528 842 1532
rect 862 1518 866 1522
rect 798 1508 802 1512
rect 850 1503 854 1507
rect 857 1503 861 1507
rect 790 1488 794 1492
rect 838 1488 842 1492
rect 766 1478 770 1482
rect 910 1728 914 1732
rect 902 1718 906 1722
rect 926 1718 930 1722
rect 918 1688 922 1692
rect 950 1738 954 1742
rect 942 1728 946 1732
rect 998 1728 1002 1732
rect 966 1718 970 1722
rect 990 1718 994 1722
rect 950 1708 954 1712
rect 942 1688 946 1692
rect 1030 1858 1034 1862
rect 1054 1868 1058 1872
rect 1110 1958 1114 1962
rect 1126 1958 1130 1962
rect 1078 1948 1082 1952
rect 1094 1948 1098 1952
rect 1142 1948 1146 1952
rect 1118 1938 1122 1942
rect 1118 1928 1122 1932
rect 1046 1848 1050 1852
rect 1038 1748 1042 1752
rect 1054 1738 1058 1742
rect 1038 1728 1042 1732
rect 1030 1718 1034 1722
rect 1022 1688 1026 1692
rect 926 1678 930 1682
rect 934 1678 938 1682
rect 1078 1888 1082 1892
rect 1094 1868 1098 1872
rect 1078 1858 1082 1862
rect 1174 2038 1178 2042
rect 1206 2048 1210 2052
rect 1198 2038 1202 2042
rect 1158 1998 1162 2002
rect 1182 1998 1186 2002
rect 1166 1978 1170 1982
rect 1190 1968 1194 1972
rect 1158 1958 1162 1962
rect 1198 1958 1202 1962
rect 1150 1928 1154 1932
rect 1254 2138 1258 2142
rect 1362 2203 1366 2207
rect 1369 2203 1373 2207
rect 1406 2288 1410 2292
rect 1414 2288 1418 2292
rect 1430 2288 1434 2292
rect 1470 2288 1474 2292
rect 1422 2268 1426 2272
rect 1502 2278 1506 2282
rect 1454 2268 1458 2272
rect 1494 2268 1498 2272
rect 1518 2268 1522 2272
rect 1438 2188 1442 2192
rect 1438 2168 1442 2172
rect 1310 2148 1314 2152
rect 1310 2128 1314 2132
rect 1294 2118 1298 2122
rect 1278 2108 1282 2112
rect 1390 2118 1394 2122
rect 1334 2068 1338 2072
rect 1358 2068 1362 2072
rect 1254 2058 1258 2062
rect 1238 2028 1242 2032
rect 1294 2018 1298 2022
rect 1254 2008 1258 2012
rect 1230 1968 1234 1972
rect 1326 1948 1330 1952
rect 1182 1938 1186 1942
rect 1222 1938 1226 1942
rect 1174 1928 1178 1932
rect 1206 1908 1210 1912
rect 1230 1928 1234 1932
rect 1214 1888 1218 1892
rect 1222 1888 1226 1892
rect 1190 1878 1194 1882
rect 1142 1868 1146 1872
rect 1222 1858 1226 1862
rect 1110 1848 1114 1852
rect 1102 1828 1106 1832
rect 1078 1808 1082 1812
rect 1094 1728 1098 1732
rect 1046 1718 1050 1722
rect 1070 1718 1074 1722
rect 902 1658 906 1662
rect 934 1658 938 1662
rect 998 1658 1002 1662
rect 1030 1658 1034 1662
rect 958 1598 962 1602
rect 918 1588 922 1592
rect 950 1588 954 1592
rect 894 1558 898 1562
rect 982 1648 986 1652
rect 1006 1648 1010 1652
rect 982 1598 986 1602
rect 998 1598 1002 1602
rect 982 1568 986 1572
rect 1022 1578 1026 1582
rect 878 1538 882 1542
rect 886 1538 890 1542
rect 902 1528 906 1532
rect 894 1518 898 1522
rect 878 1508 882 1512
rect 798 1468 802 1472
rect 814 1468 818 1472
rect 854 1468 858 1472
rect 838 1458 842 1462
rect 846 1448 850 1452
rect 806 1438 810 1442
rect 758 1428 762 1432
rect 750 1398 754 1402
rect 686 1358 690 1362
rect 710 1358 714 1362
rect 822 1438 826 1442
rect 854 1438 858 1442
rect 814 1428 818 1432
rect 798 1408 802 1412
rect 790 1368 794 1372
rect 798 1368 802 1372
rect 854 1408 858 1412
rect 870 1388 874 1392
rect 894 1378 898 1382
rect 830 1358 834 1362
rect 686 1348 690 1352
rect 758 1348 762 1352
rect 670 1338 674 1342
rect 774 1338 778 1342
rect 686 1328 690 1332
rect 694 1298 698 1302
rect 702 1278 706 1282
rect 614 1238 618 1242
rect 742 1258 746 1262
rect 742 1218 746 1222
rect 686 1188 690 1192
rect 606 1148 610 1152
rect 590 1128 594 1132
rect 710 1128 714 1132
rect 614 1108 618 1112
rect 822 1348 826 1352
rect 798 1318 802 1322
rect 782 1288 786 1292
rect 790 1268 794 1272
rect 774 1238 778 1242
rect 822 1338 826 1342
rect 990 1538 994 1542
rect 958 1528 962 1532
rect 974 1528 978 1532
rect 918 1518 922 1522
rect 926 1518 930 1522
rect 934 1458 938 1462
rect 966 1498 970 1502
rect 966 1478 970 1482
rect 1014 1518 1018 1522
rect 1014 1508 1018 1512
rect 1006 1488 1010 1492
rect 990 1478 994 1482
rect 1006 1478 1010 1482
rect 1182 1848 1186 1852
rect 1142 1828 1146 1832
rect 1158 1818 1162 1822
rect 1230 1748 1234 1752
rect 1214 1738 1218 1742
rect 1158 1728 1162 1732
rect 1174 1718 1178 1722
rect 1206 1708 1210 1712
rect 1054 1688 1058 1692
rect 1070 1688 1074 1692
rect 1110 1688 1114 1692
rect 1198 1688 1202 1692
rect 1118 1678 1122 1682
rect 1182 1678 1186 1682
rect 1094 1658 1098 1662
rect 1110 1658 1114 1662
rect 1142 1658 1146 1662
rect 1158 1638 1162 1642
rect 1206 1658 1210 1662
rect 1126 1628 1130 1632
rect 1174 1628 1178 1632
rect 1190 1628 1194 1632
rect 1110 1608 1114 1612
rect 1046 1558 1050 1562
rect 1054 1558 1058 1562
rect 1078 1558 1082 1562
rect 1038 1548 1042 1552
rect 1134 1618 1138 1622
rect 1174 1618 1178 1622
rect 1158 1598 1162 1602
rect 1246 1858 1250 1862
rect 1318 1918 1322 1922
rect 1294 1878 1298 1882
rect 1278 1868 1282 1872
rect 1270 1838 1274 1842
rect 1406 2088 1410 2092
rect 1362 2003 1366 2007
rect 1369 2003 1373 2007
rect 1350 1988 1354 1992
rect 1398 1948 1402 1952
rect 1422 2098 1426 2102
rect 1422 2088 1426 2092
rect 1422 2018 1426 2022
rect 1414 1988 1418 1992
rect 1526 2248 1530 2252
rect 1478 2228 1482 2232
rect 1518 2198 1522 2202
rect 1446 2158 1450 2162
rect 1470 2158 1474 2162
rect 1462 2148 1466 2152
rect 1454 2138 1458 2142
rect 1446 2128 1450 2132
rect 1494 2148 1498 2152
rect 1510 2138 1514 2142
rect 1494 2128 1498 2132
rect 1486 2118 1490 2122
rect 1462 2078 1466 2082
rect 1446 2068 1450 2072
rect 1462 2068 1466 2072
rect 1470 2058 1474 2062
rect 1438 2008 1442 2012
rect 1430 1998 1434 2002
rect 1454 2048 1458 2052
rect 1470 2038 1474 2042
rect 1510 2108 1514 2112
rect 1518 2108 1522 2112
rect 1494 2098 1498 2102
rect 1486 2078 1490 2082
rect 1534 2088 1538 2092
rect 1502 2068 1506 2072
rect 1510 2038 1514 2042
rect 1566 2358 1570 2362
rect 1566 2348 1570 2352
rect 1646 2518 1650 2522
rect 1662 2508 1666 2512
rect 1646 2498 1650 2502
rect 1630 2488 1634 2492
rect 1646 2468 1650 2472
rect 1678 2498 1682 2502
rect 1598 2358 1602 2362
rect 1630 2348 1634 2352
rect 1574 2338 1578 2342
rect 1582 2328 1586 2332
rect 1726 2488 1730 2492
rect 1750 2488 1754 2492
rect 1806 2648 1810 2652
rect 1822 2648 1826 2652
rect 1838 2648 1842 2652
rect 1814 2628 1818 2632
rect 1862 2608 1866 2612
rect 1798 2588 1802 2592
rect 1806 2568 1810 2572
rect 1790 2558 1794 2562
rect 1838 2558 1842 2562
rect 1806 2548 1810 2552
rect 1814 2548 1818 2552
rect 1798 2538 1802 2542
rect 1782 2518 1786 2522
rect 1790 2508 1794 2512
rect 1766 2498 1770 2502
rect 1686 2478 1690 2482
rect 1694 2478 1698 2482
rect 1726 2468 1730 2472
rect 1758 2468 1762 2472
rect 1710 2448 1714 2452
rect 1702 2438 1706 2442
rect 1742 2408 1746 2412
rect 1734 2388 1738 2392
rect 1718 2378 1722 2382
rect 1694 2358 1698 2362
rect 1662 2348 1666 2352
rect 1846 2518 1850 2522
rect 1838 2508 1842 2512
rect 1814 2488 1818 2492
rect 1830 2468 1834 2472
rect 1798 2458 1802 2462
rect 1806 2408 1810 2412
rect 1822 2428 1826 2432
rect 1822 2408 1826 2412
rect 1798 2398 1802 2402
rect 1790 2378 1794 2382
rect 1774 2358 1778 2362
rect 1790 2358 1794 2362
rect 1814 2358 1818 2362
rect 1862 2488 1866 2492
rect 1942 3128 1946 3132
rect 1942 3118 1946 3122
rect 1982 3118 1986 3122
rect 1990 3118 1994 3122
rect 1934 3108 1938 3112
rect 1934 3078 1938 3082
rect 1926 3048 1930 3052
rect 1926 3018 1930 3022
rect 1982 3098 1986 3102
rect 2014 3128 2018 3132
rect 2046 3148 2050 3152
rect 2070 3148 2074 3152
rect 2022 3118 2026 3122
rect 2054 3118 2058 3122
rect 2062 3118 2066 3122
rect 2190 3328 2194 3332
rect 2222 3318 2226 3322
rect 2182 3288 2186 3292
rect 2454 3408 2458 3412
rect 2386 3403 2390 3407
rect 2393 3403 2397 3407
rect 2358 3368 2362 3372
rect 2390 3358 2394 3362
rect 2542 3468 2546 3472
rect 2582 3468 2586 3472
rect 2534 3458 2538 3462
rect 2558 3458 2562 3462
rect 2574 3458 2578 3462
rect 2526 3448 2530 3452
rect 2542 3448 2546 3452
rect 2526 3418 2530 3422
rect 2526 3378 2530 3382
rect 2366 3348 2370 3352
rect 2486 3348 2490 3352
rect 2310 3328 2314 3332
rect 2382 3318 2386 3322
rect 2422 3318 2426 3322
rect 2318 3308 2322 3312
rect 2294 3278 2298 3282
rect 2342 3278 2346 3282
rect 2302 3258 2306 3262
rect 2342 3258 2346 3262
rect 2286 3238 2290 3242
rect 2270 3228 2274 3232
rect 2310 3248 2314 3252
rect 2294 3208 2298 3212
rect 2310 3208 2314 3212
rect 2174 3198 2178 3202
rect 2198 3198 2202 3202
rect 2294 3198 2298 3202
rect 2294 3168 2298 3172
rect 2214 3158 2218 3162
rect 2222 3158 2226 3162
rect 2158 3148 2162 3152
rect 2118 3138 2122 3142
rect 2110 3128 2114 3132
rect 2126 3128 2130 3132
rect 2118 3108 2122 3112
rect 2118 3098 2122 3102
rect 2014 3088 2018 3092
rect 1982 3068 1986 3072
rect 2014 3068 2018 3072
rect 2038 3068 2042 3072
rect 2006 3058 2010 3062
rect 1966 3048 1970 3052
rect 1982 3048 1986 3052
rect 1958 2988 1962 2992
rect 1942 2958 1946 2962
rect 1950 2938 1954 2942
rect 1902 2758 1906 2762
rect 1894 2748 1898 2752
rect 1886 2738 1890 2742
rect 1910 2728 1914 2732
rect 1910 2718 1914 2722
rect 1902 2708 1906 2712
rect 1882 2703 1886 2707
rect 1889 2703 1893 2707
rect 1878 2668 1882 2672
rect 1894 2558 1898 2562
rect 1918 2698 1922 2702
rect 2030 3058 2034 3062
rect 2070 3058 2074 3062
rect 2174 3138 2178 3142
rect 2150 3098 2154 3102
rect 2198 3148 2202 3152
rect 2222 3148 2226 3152
rect 2214 3138 2218 3142
rect 2222 3128 2226 3132
rect 2246 3128 2250 3132
rect 2230 3118 2234 3122
rect 2246 3108 2250 3112
rect 2198 3078 2202 3082
rect 2142 3058 2146 3062
rect 2166 3058 2170 3062
rect 2182 3058 2186 3062
rect 2214 3068 2218 3072
rect 2262 3108 2266 3112
rect 2254 3098 2258 3102
rect 2334 3188 2338 3192
rect 2294 3138 2298 3142
rect 2318 3128 2322 3132
rect 2310 3108 2314 3112
rect 2318 3108 2322 3112
rect 2302 3088 2306 3092
rect 2270 3078 2274 3082
rect 2366 3268 2370 3272
rect 2406 3278 2410 3282
rect 2622 3408 2626 3412
rect 2590 3328 2594 3332
rect 2606 3328 2610 3332
rect 2446 3308 2450 3312
rect 2494 3308 2498 3312
rect 2542 3308 2546 3312
rect 2910 3558 2914 3562
rect 2854 3548 2858 3552
rect 2894 3548 2898 3552
rect 2950 3568 2954 3572
rect 2926 3548 2930 3552
rect 2806 3538 2810 3542
rect 2830 3528 2834 3532
rect 2854 3518 2858 3522
rect 2906 3503 2910 3507
rect 2913 3503 2917 3507
rect 3118 3578 3122 3582
rect 3198 3578 3202 3582
rect 3238 3578 3242 3582
rect 3174 3558 3178 3562
rect 3230 3558 3234 3562
rect 3182 3548 3186 3552
rect 3222 3548 3226 3552
rect 2974 3538 2978 3542
rect 3150 3538 3154 3542
rect 3022 3528 3026 3532
rect 3038 3518 3042 3522
rect 3150 3518 3154 3522
rect 3078 3508 3082 3512
rect 2998 3498 3002 3502
rect 2902 3488 2906 3492
rect 2886 3478 2890 3482
rect 2798 3468 2802 3472
rect 2862 3468 2866 3472
rect 2878 3468 2882 3472
rect 2934 3468 2938 3472
rect 2798 3458 2802 3462
rect 2758 3448 2762 3452
rect 2750 3428 2754 3432
rect 2662 3418 2666 3422
rect 2782 3418 2786 3422
rect 2646 3398 2650 3402
rect 2774 3368 2778 3372
rect 2678 3348 2682 3352
rect 2678 3328 2682 3332
rect 2694 3298 2698 3302
rect 2438 3278 2442 3282
rect 2502 3278 2506 3282
rect 2518 3278 2522 3282
rect 2566 3278 2570 3282
rect 2510 3268 2514 3272
rect 2598 3268 2602 3272
rect 2646 3268 2650 3272
rect 2782 3338 2786 3342
rect 2814 3438 2818 3442
rect 2846 3438 2850 3442
rect 2830 3408 2834 3412
rect 2886 3448 2890 3452
rect 2870 3438 2874 3442
rect 2878 3438 2882 3442
rect 2870 3378 2874 3382
rect 2934 3418 2938 3422
rect 2878 3358 2882 3362
rect 2886 3358 2890 3362
rect 2926 3348 2930 3352
rect 2886 3338 2890 3342
rect 2902 3338 2906 3342
rect 2798 3318 2802 3322
rect 2782 3288 2786 3292
rect 2854 3278 2858 3282
rect 2390 3258 2394 3262
rect 2414 3258 2418 3262
rect 2446 3258 2450 3262
rect 2486 3258 2490 3262
rect 2542 3258 2546 3262
rect 2574 3258 2578 3262
rect 2366 3248 2370 3252
rect 2358 3168 2362 3172
rect 2350 3158 2354 3162
rect 2374 3238 2378 3242
rect 2390 3238 2394 3242
rect 2386 3203 2390 3207
rect 2393 3203 2397 3207
rect 2390 3168 2394 3172
rect 2414 3168 2418 3172
rect 2366 3128 2370 3132
rect 2326 3078 2330 3082
rect 2270 3068 2274 3072
rect 2302 3068 2306 3072
rect 2262 3058 2266 3062
rect 2278 3058 2282 3062
rect 2038 3048 2042 3052
rect 2062 3048 2066 3052
rect 2086 3048 2090 3052
rect 2126 3048 2130 3052
rect 2230 3048 2234 3052
rect 1974 2968 1978 2972
rect 2014 2968 2018 2972
rect 2030 2968 2034 2972
rect 1982 2948 1986 2952
rect 1998 2938 2002 2942
rect 2022 2938 2026 2942
rect 1982 2868 1986 2872
rect 1982 2848 1986 2852
rect 1942 2838 1946 2842
rect 1974 2838 1978 2842
rect 1942 2818 1946 2822
rect 1934 2768 1938 2772
rect 1942 2738 1946 2742
rect 1950 2728 1954 2732
rect 2006 2928 2010 2932
rect 2030 2928 2034 2932
rect 2022 2878 2026 2882
rect 2014 2858 2018 2862
rect 1998 2818 2002 2822
rect 1990 2808 1994 2812
rect 1982 2768 1986 2772
rect 2006 2788 2010 2792
rect 2014 2758 2018 2762
rect 2022 2758 2026 2762
rect 1982 2748 1986 2752
rect 2134 3038 2138 3042
rect 2102 3028 2106 3032
rect 2126 3028 2130 3032
rect 2070 3018 2074 3022
rect 2078 3018 2082 3022
rect 2062 2998 2066 3002
rect 2054 2978 2058 2982
rect 2046 2968 2050 2972
rect 2070 2928 2074 2932
rect 2110 2998 2114 3002
rect 2094 2978 2098 2982
rect 2142 2968 2146 2972
rect 2198 2968 2202 2972
rect 2214 2968 2218 2972
rect 2126 2938 2130 2942
rect 2134 2928 2138 2932
rect 2198 2938 2202 2942
rect 2222 2938 2226 2942
rect 2158 2918 2162 2922
rect 2182 2918 2186 2922
rect 2222 2918 2226 2922
rect 2046 2908 2050 2912
rect 2062 2908 2066 2912
rect 2078 2908 2082 2912
rect 2038 2898 2042 2902
rect 2070 2898 2074 2902
rect 2118 2898 2122 2902
rect 2158 2898 2162 2902
rect 2102 2878 2106 2882
rect 2270 3038 2274 3042
rect 2270 3018 2274 3022
rect 2262 2968 2266 2972
rect 2270 2958 2274 2962
rect 2398 3158 2402 3162
rect 2470 3248 2474 3252
rect 2590 3248 2594 3252
rect 2630 3248 2634 3252
rect 2478 3238 2482 3242
rect 2494 3238 2498 3242
rect 2438 3228 2442 3232
rect 2438 3178 2442 3182
rect 2422 3148 2426 3152
rect 2454 3148 2458 3152
rect 2438 3138 2442 3142
rect 2462 3128 2466 3132
rect 2398 3098 2402 3102
rect 2422 3088 2426 3092
rect 2358 3058 2362 3062
rect 2342 3028 2346 3032
rect 2334 2998 2338 3002
rect 2366 3038 2370 3042
rect 2350 2978 2354 2982
rect 2326 2968 2330 2972
rect 2318 2958 2322 2962
rect 2350 2958 2354 2962
rect 2246 2938 2250 2942
rect 2262 2918 2266 2922
rect 2238 2878 2242 2882
rect 2102 2868 2106 2872
rect 2134 2868 2138 2872
rect 2158 2868 2162 2872
rect 2198 2868 2202 2872
rect 2230 2868 2234 2872
rect 2038 2858 2042 2862
rect 2070 2858 2074 2862
rect 2086 2858 2090 2862
rect 2094 2858 2098 2862
rect 2126 2858 2130 2862
rect 2134 2858 2138 2862
rect 2150 2858 2154 2862
rect 2174 2858 2178 2862
rect 2206 2858 2210 2862
rect 2078 2848 2082 2852
rect 2198 2838 2202 2842
rect 2166 2818 2170 2822
rect 2078 2808 2082 2812
rect 2102 2808 2106 2812
rect 2222 2808 2226 2812
rect 2054 2748 2058 2752
rect 2094 2738 2098 2742
rect 2038 2728 2042 2732
rect 2046 2728 2050 2732
rect 1974 2718 1978 2722
rect 2070 2718 2074 2722
rect 2022 2708 2026 2712
rect 2246 2858 2250 2862
rect 2254 2848 2258 2852
rect 2238 2778 2242 2782
rect 2118 2758 2122 2762
rect 2110 2698 2114 2702
rect 1942 2678 1946 2682
rect 1926 2668 1930 2672
rect 1958 2668 1962 2672
rect 1998 2668 2002 2672
rect 1942 2628 1946 2632
rect 1926 2618 1930 2622
rect 1918 2608 1922 2612
rect 1942 2608 1946 2612
rect 1910 2548 1914 2552
rect 2086 2658 2090 2662
rect 2014 2628 2018 2632
rect 2094 2608 2098 2612
rect 1958 2548 1962 2552
rect 1974 2548 1978 2552
rect 2174 2748 2178 2752
rect 2206 2728 2210 2732
rect 2134 2708 2138 2712
rect 2262 2768 2266 2772
rect 2294 2928 2298 2932
rect 2302 2928 2306 2932
rect 2286 2918 2290 2922
rect 2294 2908 2298 2912
rect 2334 2948 2338 2952
rect 2398 3068 2402 3072
rect 2438 3068 2442 3072
rect 2510 3228 2514 3232
rect 2566 3228 2570 3232
rect 2502 3188 2506 3192
rect 2510 3158 2514 3162
rect 2526 3158 2530 3162
rect 2518 3148 2522 3152
rect 2510 3128 2514 3132
rect 2486 3088 2490 3092
rect 2422 3058 2426 3062
rect 2454 3058 2458 3062
rect 2430 3048 2434 3052
rect 2382 3028 2386 3032
rect 2414 3028 2418 3032
rect 2386 3003 2390 3007
rect 2393 3003 2397 3007
rect 2374 2968 2378 2972
rect 2406 2968 2410 2972
rect 2430 2968 2434 2972
rect 2398 2958 2402 2962
rect 2382 2948 2386 2952
rect 2350 2928 2354 2932
rect 2342 2908 2346 2912
rect 2382 2938 2386 2942
rect 2382 2928 2386 2932
rect 2374 2908 2378 2912
rect 2366 2888 2370 2892
rect 2302 2868 2306 2872
rect 2342 2868 2346 2872
rect 2278 2848 2282 2852
rect 2302 2848 2306 2852
rect 2318 2848 2322 2852
rect 2286 2788 2290 2792
rect 2302 2778 2306 2782
rect 2278 2768 2282 2772
rect 2286 2768 2290 2772
rect 2318 2768 2322 2772
rect 2270 2758 2274 2762
rect 2310 2758 2314 2762
rect 2270 2748 2274 2752
rect 2294 2748 2298 2752
rect 2286 2728 2290 2732
rect 2214 2708 2218 2712
rect 2246 2708 2250 2712
rect 2158 2678 2162 2682
rect 2222 2678 2226 2682
rect 2238 2678 2242 2682
rect 2254 2678 2258 2682
rect 2134 2668 2138 2672
rect 2166 2668 2170 2672
rect 2190 2668 2194 2672
rect 2214 2668 2218 2672
rect 2230 2668 2234 2672
rect 2246 2668 2250 2672
rect 2142 2658 2146 2662
rect 2110 2648 2114 2652
rect 2118 2568 2122 2572
rect 2134 2568 2138 2572
rect 2118 2558 2122 2562
rect 2150 2558 2154 2562
rect 2142 2548 2146 2552
rect 2166 2548 2170 2552
rect 1902 2538 1906 2542
rect 1974 2538 1978 2542
rect 2102 2538 2106 2542
rect 2118 2538 2122 2542
rect 1882 2503 1886 2507
rect 1889 2503 1893 2507
rect 1926 2498 1930 2502
rect 1958 2498 1962 2502
rect 1846 2478 1850 2482
rect 1854 2478 1858 2482
rect 1894 2478 1898 2482
rect 1966 2488 1970 2492
rect 1838 2458 1842 2462
rect 1894 2458 1898 2462
rect 1926 2458 1930 2462
rect 1934 2458 1938 2462
rect 1846 2448 1850 2452
rect 1854 2448 1858 2452
rect 1950 2398 1954 2402
rect 1870 2358 1874 2362
rect 1774 2348 1778 2352
rect 1806 2348 1810 2352
rect 1814 2348 1818 2352
rect 1846 2348 1850 2352
rect 1878 2348 1882 2352
rect 1670 2338 1674 2342
rect 1694 2338 1698 2342
rect 1710 2338 1714 2342
rect 1782 2338 1786 2342
rect 1614 2328 1618 2332
rect 1638 2328 1642 2332
rect 1662 2328 1666 2332
rect 1702 2328 1706 2332
rect 1590 2298 1594 2302
rect 1734 2308 1738 2312
rect 1758 2288 1762 2292
rect 1766 2288 1770 2292
rect 1750 2278 1754 2282
rect 1566 2258 1570 2262
rect 1550 2248 1554 2252
rect 1630 2248 1634 2252
rect 1614 2218 1618 2222
rect 1566 2178 1570 2182
rect 1558 2158 1562 2162
rect 1622 2198 1626 2202
rect 1694 2248 1698 2252
rect 1726 2248 1730 2252
rect 1750 2258 1754 2262
rect 1734 2208 1738 2212
rect 1742 2208 1746 2212
rect 1646 2168 1650 2172
rect 1670 2148 1674 2152
rect 1582 2138 1586 2142
rect 1606 2138 1610 2142
rect 1614 2138 1618 2142
rect 1638 2138 1642 2142
rect 1654 2138 1658 2142
rect 1662 2138 1666 2142
rect 1550 2128 1554 2132
rect 1558 2108 1562 2112
rect 1582 2108 1586 2112
rect 1550 2028 1554 2032
rect 1494 1968 1498 1972
rect 1446 1938 1450 1942
rect 1390 1918 1394 1922
rect 1390 1898 1394 1902
rect 1334 1858 1338 1862
rect 1302 1828 1306 1832
rect 1326 1828 1330 1832
rect 1362 1803 1366 1807
rect 1369 1803 1373 1807
rect 1270 1788 1274 1792
rect 1286 1788 1290 1792
rect 1246 1778 1250 1782
rect 1422 1888 1426 1892
rect 1414 1878 1418 1882
rect 1438 1858 1442 1862
rect 1438 1848 1442 1852
rect 1406 1768 1410 1772
rect 1414 1768 1418 1772
rect 1374 1758 1378 1762
rect 1358 1738 1362 1742
rect 1238 1708 1242 1712
rect 1246 1698 1250 1702
rect 1238 1688 1242 1692
rect 1374 1728 1378 1732
rect 1318 1718 1322 1722
rect 1374 1718 1378 1722
rect 1262 1698 1266 1702
rect 1398 1698 1402 1702
rect 1358 1678 1362 1682
rect 1230 1668 1234 1672
rect 1318 1668 1322 1672
rect 1334 1668 1338 1672
rect 1166 1568 1170 1572
rect 1190 1558 1194 1562
rect 1262 1638 1266 1642
rect 1230 1608 1234 1612
rect 1230 1598 1234 1602
rect 1374 1658 1378 1662
rect 1310 1638 1314 1642
rect 1342 1638 1346 1642
rect 1286 1618 1290 1622
rect 1270 1588 1274 1592
rect 1222 1578 1226 1582
rect 1206 1568 1210 1572
rect 1030 1538 1034 1542
rect 1110 1538 1114 1542
rect 1198 1538 1202 1542
rect 1054 1528 1058 1532
rect 1102 1518 1106 1522
rect 1110 1518 1114 1522
rect 1086 1488 1090 1492
rect 1142 1508 1146 1512
rect 1150 1498 1154 1502
rect 1150 1488 1154 1492
rect 1182 1508 1186 1512
rect 1174 1488 1178 1492
rect 1190 1488 1194 1492
rect 998 1468 1002 1472
rect 1046 1468 1050 1472
rect 1070 1468 1074 1472
rect 950 1438 954 1442
rect 958 1438 962 1442
rect 958 1418 962 1422
rect 942 1398 946 1402
rect 918 1368 922 1372
rect 950 1358 954 1362
rect 910 1348 914 1352
rect 934 1338 938 1342
rect 830 1328 834 1332
rect 894 1328 898 1332
rect 814 1278 818 1282
rect 814 1258 818 1262
rect 850 1303 854 1307
rect 857 1303 861 1307
rect 918 1318 922 1322
rect 926 1318 930 1322
rect 902 1308 906 1312
rect 918 1308 922 1312
rect 926 1278 930 1282
rect 934 1218 938 1222
rect 894 1198 898 1202
rect 886 1188 890 1192
rect 846 1178 850 1182
rect 806 1138 810 1142
rect 710 1118 714 1122
rect 758 1118 762 1122
rect 614 1088 618 1092
rect 694 1088 698 1092
rect 846 1148 850 1152
rect 862 1148 866 1152
rect 878 1148 882 1152
rect 830 1128 834 1132
rect 798 1108 802 1112
rect 850 1103 854 1107
rect 857 1103 861 1107
rect 742 1098 746 1102
rect 782 1098 786 1102
rect 822 1098 826 1102
rect 838 1098 842 1102
rect 822 1088 826 1092
rect 710 1078 714 1082
rect 694 1068 698 1072
rect 550 988 554 992
rect 454 938 458 942
rect 486 938 490 942
rect 534 938 538 942
rect 446 928 450 932
rect 462 898 466 902
rect 398 888 402 892
rect 414 888 418 892
rect 454 888 458 892
rect 446 878 450 882
rect 470 878 474 882
rect 510 928 514 932
rect 502 898 506 902
rect 494 888 498 892
rect 534 918 538 922
rect 526 898 530 902
rect 526 888 530 892
rect 918 1168 922 1172
rect 902 1158 906 1162
rect 910 1148 914 1152
rect 926 1148 930 1152
rect 966 1348 970 1352
rect 982 1348 986 1352
rect 990 1348 994 1352
rect 1030 1458 1034 1462
rect 1054 1458 1058 1462
rect 1094 1468 1098 1472
rect 1142 1468 1146 1472
rect 1198 1468 1202 1472
rect 1206 1468 1210 1472
rect 1022 1368 1026 1372
rect 958 1338 962 1342
rect 990 1338 994 1342
rect 1006 1338 1010 1342
rect 966 1308 970 1312
rect 950 1268 954 1272
rect 990 1298 994 1302
rect 1006 1318 1010 1322
rect 998 1278 1002 1282
rect 974 1258 978 1262
rect 966 1148 970 1152
rect 894 1138 898 1142
rect 942 1138 946 1142
rect 942 1128 946 1132
rect 822 1068 826 1072
rect 886 1068 890 1072
rect 1086 1418 1090 1422
rect 1118 1398 1122 1402
rect 1126 1368 1130 1372
rect 1070 1348 1074 1352
rect 1134 1348 1138 1352
rect 1086 1318 1090 1322
rect 1070 1308 1074 1312
rect 1086 1308 1090 1312
rect 1030 1298 1034 1302
rect 1030 1288 1034 1292
rect 1238 1468 1242 1472
rect 1150 1458 1154 1462
rect 1182 1448 1186 1452
rect 1206 1448 1210 1452
rect 1166 1418 1170 1422
rect 1166 1398 1170 1402
rect 1166 1368 1170 1372
rect 1350 1608 1354 1612
rect 1362 1603 1366 1607
rect 1369 1603 1373 1607
rect 1326 1548 1330 1552
rect 1518 1958 1522 1962
rect 1478 1948 1482 1952
rect 1462 1928 1466 1932
rect 1510 1928 1514 1932
rect 1526 1928 1530 1932
rect 1486 1888 1490 1892
rect 1534 1898 1538 1902
rect 1526 1888 1530 1892
rect 1510 1878 1514 1882
rect 1582 2068 1586 2072
rect 1638 2068 1642 2072
rect 1566 2038 1570 2042
rect 1702 2128 1706 2132
rect 1726 2108 1730 2112
rect 1710 2088 1714 2092
rect 1718 2078 1722 2082
rect 1742 2068 1746 2072
rect 1694 2058 1698 2062
rect 1622 2038 1626 2042
rect 1654 2008 1658 2012
rect 1590 1998 1594 2002
rect 1582 1968 1586 1972
rect 1630 1968 1634 1972
rect 1742 2048 1746 2052
rect 1854 2338 1858 2342
rect 1846 2328 1850 2332
rect 1870 2318 1874 2322
rect 1902 2318 1906 2322
rect 1918 2318 1922 2322
rect 1862 2308 1866 2312
rect 1882 2303 1886 2307
rect 1889 2303 1893 2307
rect 1862 2278 1866 2282
rect 1774 2268 1778 2272
rect 1798 2268 1802 2272
rect 1822 2268 1826 2272
rect 1870 2268 1874 2272
rect 1910 2268 1914 2272
rect 1782 2248 1786 2252
rect 1758 2238 1762 2242
rect 1774 2238 1778 2242
rect 1838 2258 1842 2262
rect 1838 2248 1842 2252
rect 1814 2208 1818 2212
rect 1878 2258 1882 2262
rect 1862 2188 1866 2192
rect 1790 2178 1794 2182
rect 1766 2168 1770 2172
rect 1814 2158 1818 2162
rect 1846 2158 1850 2162
rect 1862 2158 1866 2162
rect 1774 2148 1778 2152
rect 1798 2148 1802 2152
rect 1798 2138 1802 2142
rect 1774 2098 1778 2102
rect 1766 2088 1770 2092
rect 1766 2078 1770 2082
rect 1830 2138 1834 2142
rect 1982 2518 1986 2522
rect 2014 2508 2018 2512
rect 2006 2478 2010 2482
rect 1998 2388 2002 2392
rect 1982 2358 1986 2362
rect 1958 2338 1962 2342
rect 2094 2528 2098 2532
rect 2142 2528 2146 2532
rect 2038 2508 2042 2512
rect 2054 2508 2058 2512
rect 2030 2478 2034 2482
rect 2078 2468 2082 2472
rect 2062 2458 2066 2462
rect 2086 2458 2090 2462
rect 2038 2448 2042 2452
rect 2022 2418 2026 2422
rect 2078 2438 2082 2442
rect 2038 2388 2042 2392
rect 2022 2358 2026 2362
rect 2022 2348 2026 2352
rect 2014 2338 2018 2342
rect 2038 2338 2042 2342
rect 1990 2328 1994 2332
rect 1982 2318 1986 2322
rect 1974 2308 1978 2312
rect 1990 2288 1994 2292
rect 1998 2288 2002 2292
rect 1950 2268 1954 2272
rect 1902 2248 1906 2252
rect 1926 2248 1930 2252
rect 1958 2218 1962 2222
rect 1974 2218 1978 2222
rect 1926 2188 1930 2192
rect 1966 2188 1970 2192
rect 1918 2168 1922 2172
rect 1902 2148 1906 2152
rect 1950 2168 1954 2172
rect 1958 2158 1962 2162
rect 1982 2158 1986 2162
rect 1918 2138 1922 2142
rect 1886 2128 1890 2132
rect 1846 2118 1850 2122
rect 1878 2118 1882 2122
rect 2070 2368 2074 2372
rect 2046 2328 2050 2332
rect 2038 2298 2042 2302
rect 2062 2298 2066 2302
rect 2102 2498 2106 2502
rect 2158 2498 2162 2502
rect 2142 2468 2146 2472
rect 2118 2458 2122 2462
rect 2102 2438 2106 2442
rect 2126 2438 2130 2442
rect 2014 2268 2018 2272
rect 2094 2268 2098 2272
rect 1998 2248 2002 2252
rect 2182 2538 2186 2542
rect 2182 2518 2186 2522
rect 2190 2508 2194 2512
rect 2246 2658 2250 2662
rect 2262 2648 2266 2652
rect 2318 2658 2322 2662
rect 2294 2628 2298 2632
rect 2310 2628 2314 2632
rect 2278 2618 2282 2622
rect 2206 2608 2210 2612
rect 2302 2588 2306 2592
rect 2318 2588 2322 2592
rect 2262 2578 2266 2582
rect 2342 2838 2346 2842
rect 2342 2808 2346 2812
rect 2398 2878 2402 2882
rect 2422 2948 2426 2952
rect 2430 2938 2434 2942
rect 2422 2888 2426 2892
rect 2414 2878 2418 2882
rect 2382 2858 2386 2862
rect 2386 2803 2390 2807
rect 2393 2803 2397 2807
rect 2390 2788 2394 2792
rect 2334 2758 2338 2762
rect 2366 2758 2370 2762
rect 2342 2748 2346 2752
rect 2366 2748 2370 2752
rect 2374 2738 2378 2742
rect 2366 2708 2370 2712
rect 2350 2678 2354 2682
rect 2342 2668 2346 2672
rect 2422 2868 2426 2872
rect 2446 3038 2450 3042
rect 2462 3038 2466 3042
rect 2462 3008 2466 3012
rect 2462 2978 2466 2982
rect 2478 3038 2482 3042
rect 2494 3078 2498 3082
rect 2486 3018 2490 3022
rect 2542 3148 2546 3152
rect 2566 3148 2570 3152
rect 2582 3148 2586 3152
rect 2566 3138 2570 3142
rect 2798 3258 2802 3262
rect 2622 3178 2626 3182
rect 2606 3168 2610 3172
rect 2638 3148 2642 3152
rect 2606 3138 2610 3142
rect 2598 3118 2602 3122
rect 2534 3098 2538 3102
rect 2590 3098 2594 3102
rect 2622 3098 2626 3102
rect 2630 3098 2634 3102
rect 2566 3078 2570 3082
rect 2510 3008 2514 3012
rect 2502 2978 2506 2982
rect 2694 3248 2698 3252
rect 2662 3098 2666 3102
rect 2654 3078 2658 3082
rect 2574 3068 2578 3072
rect 2566 3058 2570 3062
rect 2590 3058 2594 3062
rect 2606 3058 2610 3062
rect 2542 3038 2546 3042
rect 2566 3038 2570 3042
rect 2534 3028 2538 3032
rect 2566 2978 2570 2982
rect 2478 2968 2482 2972
rect 2526 2968 2530 2972
rect 2542 2968 2546 2972
rect 2454 2958 2458 2962
rect 2462 2958 2466 2962
rect 2470 2958 2474 2962
rect 2446 2948 2450 2952
rect 2454 2938 2458 2942
rect 2518 2948 2522 2952
rect 2454 2888 2458 2892
rect 2494 2938 2498 2942
rect 2486 2918 2490 2922
rect 2534 2918 2538 2922
rect 2542 2898 2546 2902
rect 2574 2938 2578 2942
rect 2670 3078 2674 3082
rect 2686 3108 2690 3112
rect 2742 3198 2746 3202
rect 2758 3198 2762 3202
rect 2702 3108 2706 3112
rect 2670 3058 2674 3062
rect 2774 3138 2778 3142
rect 2758 3128 2762 3132
rect 2894 3328 2898 3332
rect 2870 3308 2874 3312
rect 2906 3303 2910 3307
rect 2913 3303 2917 3307
rect 2894 3288 2898 3292
rect 2918 3278 2922 3282
rect 3038 3488 3042 3492
rect 3014 3458 3018 3462
rect 3118 3488 3122 3492
rect 3158 3508 3162 3512
rect 3190 3508 3194 3512
rect 3158 3498 3162 3502
rect 3118 3478 3122 3482
rect 2966 3448 2970 3452
rect 3006 3448 3010 3452
rect 2974 3438 2978 3442
rect 2982 3438 2986 3442
rect 3030 3438 3034 3442
rect 2950 3398 2954 3402
rect 2958 3388 2962 3392
rect 2950 3378 2954 3382
rect 2966 3358 2970 3362
rect 2966 3338 2970 3342
rect 2990 3408 2994 3412
rect 2982 3388 2986 3392
rect 2974 3328 2978 3332
rect 2926 3268 2930 3272
rect 2918 3248 2922 3252
rect 2862 3168 2866 3172
rect 2926 3168 2930 3172
rect 2950 3308 2954 3312
rect 2982 3308 2986 3312
rect 3006 3378 3010 3382
rect 3022 3378 3026 3382
rect 2998 3358 3002 3362
rect 3014 3348 3018 3352
rect 2998 3338 3002 3342
rect 3030 3308 3034 3312
rect 3014 3298 3018 3302
rect 3014 3278 3018 3282
rect 2950 3268 2954 3272
rect 2974 3268 2978 3272
rect 3014 3268 3018 3272
rect 2958 3258 2962 3262
rect 2982 3258 2986 3262
rect 3070 3458 3074 3462
rect 3110 3458 3114 3462
rect 3134 3448 3138 3452
rect 3142 3438 3146 3442
rect 3062 3418 3066 3422
rect 3166 3418 3170 3422
rect 3174 3418 3178 3422
rect 3094 3368 3098 3372
rect 3054 3358 3058 3362
rect 3110 3338 3114 3342
rect 3046 3318 3050 3322
rect 3062 3318 3066 3322
rect 3038 3298 3042 3302
rect 3038 3278 3042 3282
rect 3022 3258 3026 3262
rect 3102 3318 3106 3322
rect 3086 3308 3090 3312
rect 3070 3298 3074 3302
rect 3054 3258 3058 3262
rect 3062 3248 3066 3252
rect 3038 3238 3042 3242
rect 3054 3188 3058 3192
rect 3014 3148 3018 3152
rect 3094 3278 3098 3282
rect 3086 3268 3090 3272
rect 3078 3218 3082 3222
rect 3078 3158 3082 3162
rect 3214 3538 3218 3542
rect 3214 3488 3218 3492
rect 3214 3448 3218 3452
rect 3230 3448 3234 3452
rect 3318 3568 3322 3572
rect 3342 3568 3346 3572
rect 3454 3568 3458 3572
rect 3478 3568 3482 3572
rect 3678 3568 3682 3572
rect 3686 3568 3690 3572
rect 3246 3548 3250 3552
rect 3278 3548 3282 3552
rect 3286 3548 3290 3552
rect 3326 3548 3330 3552
rect 3254 3528 3258 3532
rect 3262 3508 3266 3512
rect 3310 3538 3314 3542
rect 3294 3518 3298 3522
rect 3294 3508 3298 3512
rect 3278 3498 3282 3502
rect 3334 3518 3338 3522
rect 3438 3558 3442 3562
rect 3350 3548 3354 3552
rect 3374 3548 3378 3552
rect 3390 3548 3394 3552
rect 3430 3548 3434 3552
rect 3350 3518 3354 3522
rect 3310 3498 3314 3502
rect 3302 3478 3306 3482
rect 3358 3468 3362 3472
rect 3270 3448 3274 3452
rect 3286 3448 3290 3452
rect 3238 3438 3242 3442
rect 3254 3438 3258 3442
rect 3246 3418 3250 3422
rect 3254 3418 3258 3422
rect 3270 3418 3274 3422
rect 3286 3418 3290 3422
rect 3222 3408 3226 3412
rect 3198 3388 3202 3392
rect 3190 3378 3194 3382
rect 3246 3388 3250 3392
rect 3278 3378 3282 3382
rect 3190 3368 3194 3372
rect 3222 3368 3226 3372
rect 3246 3368 3250 3372
rect 3254 3368 3258 3372
rect 3126 3348 3130 3352
rect 3166 3348 3170 3352
rect 3134 3338 3138 3342
rect 3118 3288 3122 3292
rect 3150 3288 3154 3292
rect 3206 3358 3210 3362
rect 3230 3358 3234 3362
rect 3270 3358 3274 3362
rect 3206 3328 3210 3332
rect 3174 3308 3178 3312
rect 3166 3278 3170 3282
rect 3158 3268 3162 3272
rect 3182 3278 3186 3282
rect 3278 3348 3282 3352
rect 3246 3338 3250 3342
rect 3270 3328 3274 3332
rect 3262 3308 3266 3312
rect 3278 3308 3282 3312
rect 3246 3298 3250 3302
rect 3230 3288 3234 3292
rect 3246 3288 3250 3292
rect 3238 3278 3242 3282
rect 3246 3278 3250 3282
rect 3222 3268 3226 3272
rect 3126 3258 3130 3262
rect 3174 3258 3178 3262
rect 3102 3248 3106 3252
rect 2998 3138 3002 3142
rect 3094 3128 3098 3132
rect 2934 3118 2938 3122
rect 2990 3118 2994 3122
rect 3110 3118 3114 3122
rect 2862 3088 2866 3092
rect 2854 3078 2858 3082
rect 2806 3068 2810 3072
rect 2694 3058 2698 3062
rect 2710 3058 2714 3062
rect 2758 3058 2762 3062
rect 2678 3048 2682 3052
rect 2646 3038 2650 3042
rect 2694 3038 2698 3042
rect 2622 2978 2626 2982
rect 2822 3028 2826 3032
rect 2726 2998 2730 3002
rect 2750 2998 2754 3002
rect 2718 2978 2722 2982
rect 2678 2948 2682 2952
rect 2906 3103 2910 3107
rect 2913 3103 2917 3107
rect 2974 3078 2978 3082
rect 2878 3048 2882 3052
rect 2878 3018 2882 3022
rect 2662 2938 2666 2942
rect 2742 2938 2746 2942
rect 2766 2938 2770 2942
rect 2622 2928 2626 2932
rect 2614 2918 2618 2922
rect 2606 2908 2610 2912
rect 2662 2908 2666 2912
rect 2686 2908 2690 2912
rect 2630 2878 2634 2882
rect 2646 2878 2650 2882
rect 2758 2918 2762 2922
rect 2766 2888 2770 2892
rect 2854 2938 2858 2942
rect 3022 3008 3026 3012
rect 2982 2968 2986 2972
rect 2958 2958 2962 2962
rect 2926 2948 2930 2952
rect 2870 2918 2874 2922
rect 2918 2918 2922 2922
rect 2798 2908 2802 2912
rect 2906 2903 2910 2907
rect 2913 2903 2917 2907
rect 2902 2888 2906 2892
rect 2814 2878 2818 2882
rect 2830 2878 2834 2882
rect 2614 2868 2618 2872
rect 2694 2868 2698 2872
rect 2750 2868 2754 2872
rect 2758 2868 2762 2872
rect 2462 2828 2466 2832
rect 2446 2818 2450 2822
rect 2438 2808 2442 2812
rect 2574 2858 2578 2862
rect 2630 2858 2634 2862
rect 2662 2858 2666 2862
rect 2518 2848 2522 2852
rect 2542 2848 2546 2852
rect 2590 2848 2594 2852
rect 2598 2848 2602 2852
rect 2622 2848 2626 2852
rect 2646 2848 2650 2852
rect 2502 2838 2506 2842
rect 2518 2818 2522 2822
rect 2534 2808 2538 2812
rect 2478 2788 2482 2792
rect 2478 2758 2482 2762
rect 2398 2728 2402 2732
rect 2422 2738 2426 2742
rect 2446 2738 2450 2742
rect 2454 2728 2458 2732
rect 2438 2718 2442 2722
rect 2462 2698 2466 2702
rect 2446 2688 2450 2692
rect 2414 2678 2418 2682
rect 2366 2668 2370 2672
rect 2446 2668 2450 2672
rect 2414 2658 2418 2662
rect 2382 2648 2386 2652
rect 2414 2648 2418 2652
rect 2446 2648 2450 2652
rect 2406 2628 2410 2632
rect 2374 2608 2378 2612
rect 2386 2603 2390 2607
rect 2393 2603 2397 2607
rect 2406 2598 2410 2602
rect 2390 2578 2394 2582
rect 2422 2568 2426 2572
rect 2542 2748 2546 2752
rect 2558 2728 2562 2732
rect 2646 2818 2650 2822
rect 2630 2768 2634 2772
rect 2606 2758 2610 2762
rect 2686 2848 2690 2852
rect 2710 2848 2714 2852
rect 2718 2838 2722 2842
rect 2694 2828 2698 2832
rect 2678 2798 2682 2802
rect 2662 2758 2666 2762
rect 2598 2718 2602 2722
rect 2542 2668 2546 2672
rect 2502 2638 2506 2642
rect 2374 2558 2378 2562
rect 2382 2558 2386 2562
rect 2454 2558 2458 2562
rect 2494 2558 2498 2562
rect 2326 2548 2330 2552
rect 2342 2538 2346 2542
rect 2262 2528 2266 2532
rect 2302 2528 2306 2532
rect 2318 2528 2322 2532
rect 2334 2528 2338 2532
rect 2246 2518 2250 2522
rect 2230 2508 2234 2512
rect 2206 2488 2210 2492
rect 2238 2488 2242 2492
rect 2286 2488 2290 2492
rect 2310 2488 2314 2492
rect 2198 2468 2202 2472
rect 2222 2458 2226 2462
rect 2182 2438 2186 2442
rect 2190 2428 2194 2432
rect 2302 2468 2306 2472
rect 2334 2518 2338 2522
rect 2350 2458 2354 2462
rect 2286 2438 2290 2442
rect 2246 2428 2250 2432
rect 2222 2418 2226 2422
rect 2278 2418 2282 2422
rect 2262 2408 2266 2412
rect 2430 2548 2434 2552
rect 2406 2528 2410 2532
rect 2390 2518 2394 2522
rect 2382 2508 2386 2512
rect 2422 2518 2426 2522
rect 2438 2518 2442 2522
rect 2406 2498 2410 2502
rect 2374 2488 2378 2492
rect 2430 2498 2434 2502
rect 2470 2498 2474 2502
rect 2366 2468 2370 2472
rect 2366 2448 2370 2452
rect 2358 2408 2362 2412
rect 2278 2398 2282 2402
rect 2166 2388 2170 2392
rect 2294 2378 2298 2382
rect 2302 2358 2306 2362
rect 2254 2348 2258 2352
rect 2286 2348 2290 2352
rect 2158 2338 2162 2342
rect 2158 2318 2162 2322
rect 2174 2318 2178 2322
rect 2126 2268 2130 2272
rect 2166 2268 2170 2272
rect 2310 2338 2314 2342
rect 2326 2338 2330 2342
rect 2334 2328 2338 2332
rect 2390 2458 2394 2462
rect 2422 2448 2426 2452
rect 2446 2458 2450 2462
rect 2734 2788 2738 2792
rect 2726 2768 2730 2772
rect 2742 2758 2746 2762
rect 2710 2748 2714 2752
rect 2646 2738 2650 2742
rect 2662 2738 2666 2742
rect 2686 2738 2690 2742
rect 2638 2718 2642 2722
rect 2654 2718 2658 2722
rect 2630 2698 2634 2702
rect 2646 2698 2650 2702
rect 2678 2698 2682 2702
rect 2638 2688 2642 2692
rect 2734 2728 2738 2732
rect 2702 2708 2706 2712
rect 2678 2668 2682 2672
rect 2702 2668 2706 2672
rect 2598 2658 2602 2662
rect 2558 2628 2562 2632
rect 2542 2608 2546 2612
rect 2534 2598 2538 2602
rect 2510 2558 2514 2562
rect 2534 2558 2538 2562
rect 2510 2538 2514 2542
rect 2550 2568 2554 2572
rect 2582 2568 2586 2572
rect 2654 2648 2658 2652
rect 2662 2648 2666 2652
rect 2718 2648 2722 2652
rect 2670 2638 2674 2642
rect 2742 2638 2746 2642
rect 2782 2858 2786 2862
rect 2814 2858 2818 2862
rect 2774 2788 2778 2792
rect 2918 2808 2922 2812
rect 2934 2808 2938 2812
rect 2918 2788 2922 2792
rect 2790 2768 2794 2772
rect 2862 2758 2866 2762
rect 2782 2748 2786 2752
rect 2766 2738 2770 2742
rect 2790 2738 2794 2742
rect 2822 2738 2826 2742
rect 2774 2728 2778 2732
rect 2774 2698 2778 2702
rect 2798 2668 2802 2672
rect 2854 2748 2858 2752
rect 2878 2748 2882 2752
rect 2918 2748 2922 2752
rect 2846 2738 2850 2742
rect 2830 2728 2834 2732
rect 2814 2668 2818 2672
rect 2758 2638 2762 2642
rect 2774 2628 2778 2632
rect 2670 2598 2674 2602
rect 2798 2638 2802 2642
rect 2806 2628 2810 2632
rect 2822 2638 2826 2642
rect 2862 2698 2866 2702
rect 2854 2668 2858 2672
rect 2846 2648 2850 2652
rect 2838 2588 2842 2592
rect 2702 2578 2706 2582
rect 2782 2578 2786 2582
rect 2814 2578 2818 2582
rect 2830 2578 2834 2582
rect 2838 2578 2842 2582
rect 2830 2568 2834 2572
rect 2718 2558 2722 2562
rect 2790 2558 2794 2562
rect 2542 2518 2546 2522
rect 2534 2508 2538 2512
rect 2550 2508 2554 2512
rect 2494 2478 2498 2482
rect 2478 2448 2482 2452
rect 2438 2438 2442 2442
rect 2386 2403 2390 2407
rect 2393 2403 2397 2407
rect 2470 2398 2474 2402
rect 2422 2348 2426 2352
rect 2486 2348 2490 2352
rect 2382 2338 2386 2342
rect 2438 2338 2442 2342
rect 2422 2328 2426 2332
rect 2262 2288 2266 2292
rect 2326 2288 2330 2292
rect 2366 2288 2370 2292
rect 2374 2288 2378 2292
rect 2118 2258 2122 2262
rect 2030 2248 2034 2252
rect 2022 2238 2026 2242
rect 2006 2228 2010 2232
rect 2046 2228 2050 2232
rect 2014 2218 2018 2222
rect 2006 2208 2010 2212
rect 2102 2248 2106 2252
rect 2158 2198 2162 2202
rect 1998 2188 2002 2192
rect 1958 2148 1962 2152
rect 1966 2148 1970 2152
rect 1966 2128 1970 2132
rect 1942 2108 1946 2112
rect 1882 2103 1886 2107
rect 1889 2103 1893 2107
rect 1870 2098 1874 2102
rect 1806 2078 1810 2082
rect 1830 2078 1834 2082
rect 1870 2078 1874 2082
rect 1894 2078 1898 2082
rect 2054 2178 2058 2182
rect 2502 2438 2506 2442
rect 2534 2398 2538 2402
rect 2518 2378 2522 2382
rect 2510 2368 2514 2372
rect 2582 2548 2586 2552
rect 2598 2548 2602 2552
rect 2654 2548 2658 2552
rect 2662 2548 2666 2552
rect 2686 2548 2690 2552
rect 2710 2548 2714 2552
rect 2574 2528 2578 2532
rect 2638 2528 2642 2532
rect 2630 2518 2634 2522
rect 2566 2498 2570 2502
rect 2606 2498 2610 2502
rect 2630 2498 2634 2502
rect 2742 2538 2746 2542
rect 2750 2538 2754 2542
rect 2774 2538 2778 2542
rect 2806 2538 2810 2542
rect 2686 2488 2690 2492
rect 2726 2498 2730 2502
rect 2798 2528 2802 2532
rect 2766 2508 2770 2512
rect 2710 2478 2714 2482
rect 2614 2468 2618 2472
rect 2694 2468 2698 2472
rect 2734 2468 2738 2472
rect 2750 2468 2754 2472
rect 2710 2458 2714 2462
rect 2558 2378 2562 2382
rect 2550 2358 2554 2362
rect 2566 2368 2570 2372
rect 2534 2338 2538 2342
rect 2614 2368 2618 2372
rect 2606 2358 2610 2362
rect 2574 2348 2578 2352
rect 2590 2348 2594 2352
rect 2590 2328 2594 2332
rect 2598 2328 2602 2332
rect 2518 2308 2522 2312
rect 2582 2298 2586 2302
rect 2502 2288 2506 2292
rect 2358 2278 2362 2282
rect 2414 2278 2418 2282
rect 2422 2278 2426 2282
rect 2462 2278 2466 2282
rect 2382 2268 2386 2272
rect 2518 2278 2522 2282
rect 2654 2358 2658 2362
rect 2630 2338 2634 2342
rect 2662 2338 2666 2342
rect 2654 2288 2658 2292
rect 2646 2278 2650 2282
rect 2446 2268 2450 2272
rect 2486 2268 2490 2272
rect 2494 2268 2498 2272
rect 2558 2268 2562 2272
rect 2590 2268 2594 2272
rect 2622 2268 2626 2272
rect 2638 2268 2642 2272
rect 2358 2258 2362 2262
rect 2358 2248 2362 2252
rect 2406 2248 2410 2252
rect 2158 2178 2162 2182
rect 2222 2178 2226 2182
rect 2278 2168 2282 2172
rect 2182 2158 2186 2162
rect 2238 2158 2242 2162
rect 2206 2148 2210 2152
rect 2094 2138 2098 2142
rect 1974 2098 1978 2102
rect 1990 2098 1994 2102
rect 1790 2068 1794 2072
rect 1798 2068 1802 2072
rect 1766 2048 1770 2052
rect 1782 2048 1786 2052
rect 1806 2048 1810 2052
rect 1822 2048 1826 2052
rect 1774 2038 1778 2042
rect 1830 2038 1834 2042
rect 1750 2028 1754 2032
rect 1790 2028 1794 2032
rect 1758 1978 1762 1982
rect 1710 1968 1714 1972
rect 1742 1968 1746 1972
rect 1782 1978 1786 1982
rect 1606 1958 1610 1962
rect 1758 1958 1762 1962
rect 1598 1948 1602 1952
rect 1662 1948 1666 1952
rect 1718 1948 1722 1952
rect 1566 1938 1570 1942
rect 1590 1938 1594 1942
rect 1558 1928 1562 1932
rect 1558 1908 1562 1912
rect 1574 1898 1578 1902
rect 1550 1878 1554 1882
rect 1526 1868 1530 1872
rect 1590 1868 1594 1872
rect 1478 1858 1482 1862
rect 1518 1858 1522 1862
rect 1526 1838 1530 1842
rect 1534 1838 1538 1842
rect 1454 1778 1458 1782
rect 1454 1768 1458 1772
rect 1478 1768 1482 1772
rect 1446 1758 1450 1762
rect 1494 1758 1498 1762
rect 1614 1938 1618 1942
rect 1630 1938 1634 1942
rect 1622 1928 1626 1932
rect 1862 2068 1866 2072
rect 1870 2068 1874 2072
rect 1886 2068 1890 2072
rect 1934 2068 1938 2072
rect 1854 2028 1858 2032
rect 1918 2058 1922 2062
rect 1942 2058 1946 2062
rect 1902 2048 1906 2052
rect 1926 2028 1930 2032
rect 1958 2028 1962 2032
rect 1870 1978 1874 1982
rect 1838 1968 1842 1972
rect 1814 1958 1818 1962
rect 1830 1958 1834 1962
rect 1822 1948 1826 1952
rect 1726 1938 1730 1942
rect 1782 1938 1786 1942
rect 1718 1928 1722 1932
rect 1694 1918 1698 1922
rect 1718 1918 1722 1922
rect 1686 1908 1690 1912
rect 1694 1908 1698 1912
rect 1646 1898 1650 1902
rect 1678 1898 1682 1902
rect 1854 1958 1858 1962
rect 1846 1938 1850 1942
rect 1790 1908 1794 1912
rect 1822 1908 1826 1912
rect 1750 1898 1754 1902
rect 1790 1898 1794 1902
rect 1622 1888 1626 1892
rect 1670 1878 1674 1882
rect 1806 1878 1810 1882
rect 1566 1838 1570 1842
rect 1574 1838 1578 1842
rect 1550 1798 1554 1802
rect 1566 1758 1570 1762
rect 1598 1828 1602 1832
rect 1614 1848 1618 1852
rect 1582 1778 1586 1782
rect 1598 1778 1602 1782
rect 1606 1778 1610 1782
rect 1606 1758 1610 1762
rect 1494 1738 1498 1742
rect 1454 1728 1458 1732
rect 1422 1688 1426 1692
rect 1414 1668 1418 1672
rect 1510 1718 1514 1722
rect 1486 1708 1490 1712
rect 1470 1698 1474 1702
rect 1462 1678 1466 1682
rect 1430 1668 1434 1672
rect 1470 1668 1474 1672
rect 1478 1668 1482 1672
rect 1526 1728 1530 1732
rect 1502 1668 1506 1672
rect 1518 1698 1522 1702
rect 1526 1678 1530 1682
rect 1558 1748 1562 1752
rect 1590 1748 1594 1752
rect 1494 1638 1498 1642
rect 1470 1628 1474 1632
rect 1454 1578 1458 1582
rect 1462 1578 1466 1582
rect 1438 1568 1442 1572
rect 1550 1608 1554 1612
rect 1518 1568 1522 1572
rect 1406 1558 1410 1562
rect 1502 1558 1506 1562
rect 1678 1868 1682 1872
rect 1622 1798 1626 1802
rect 1622 1748 1626 1752
rect 1566 1738 1570 1742
rect 1622 1738 1626 1742
rect 1662 1848 1666 1852
rect 1646 1828 1650 1832
rect 1638 1768 1642 1772
rect 1646 1758 1650 1762
rect 1638 1738 1642 1742
rect 1630 1708 1634 1712
rect 1606 1698 1610 1702
rect 1622 1698 1626 1702
rect 1862 1938 1866 1942
rect 2070 2078 2074 2082
rect 1990 1968 1994 1972
rect 2022 1988 2026 1992
rect 2030 1978 2034 1982
rect 2014 1958 2018 1962
rect 2022 1958 2026 1962
rect 1966 1948 1970 1952
rect 1982 1938 1986 1942
rect 1918 1928 1922 1932
rect 2150 2048 2154 2052
rect 2110 2038 2114 2042
rect 2142 2008 2146 2012
rect 2206 2128 2210 2132
rect 2190 2108 2194 2112
rect 2326 2218 2330 2222
rect 2302 2188 2306 2192
rect 2318 2188 2322 2192
rect 2294 2158 2298 2162
rect 2246 2138 2250 2142
rect 2222 2128 2226 2132
rect 2222 2088 2226 2092
rect 2238 2088 2242 2092
rect 2214 2078 2218 2082
rect 2166 2068 2170 2072
rect 2222 2068 2226 2072
rect 2222 2058 2226 2062
rect 2174 2048 2178 2052
rect 2190 1958 2194 1962
rect 2126 1948 2130 1952
rect 2222 2048 2226 2052
rect 2254 2128 2258 2132
rect 2270 2098 2274 2102
rect 2310 2138 2314 2142
rect 2302 2088 2306 2092
rect 2342 2208 2346 2212
rect 2350 2208 2354 2212
rect 2386 2203 2390 2207
rect 2393 2203 2397 2207
rect 2374 2198 2378 2202
rect 2438 2238 2442 2242
rect 2550 2258 2554 2262
rect 2582 2258 2586 2262
rect 2486 2248 2490 2252
rect 2614 2258 2618 2262
rect 2630 2258 2634 2262
rect 2470 2238 2474 2242
rect 2454 2208 2458 2212
rect 2430 2188 2434 2192
rect 2494 2238 2498 2242
rect 2518 2188 2522 2192
rect 2462 2178 2466 2182
rect 2470 2178 2474 2182
rect 2486 2178 2490 2182
rect 2374 2168 2378 2172
rect 2462 2158 2466 2162
rect 2342 2138 2346 2142
rect 2334 2098 2338 2102
rect 2358 2138 2362 2142
rect 2390 2138 2394 2142
rect 2430 2138 2434 2142
rect 2366 2128 2370 2132
rect 2454 2138 2458 2142
rect 2446 2128 2450 2132
rect 2422 2108 2426 2112
rect 2350 2088 2354 2092
rect 2358 2088 2362 2092
rect 2398 2088 2402 2092
rect 2414 2088 2418 2092
rect 2294 2078 2298 2082
rect 2302 2078 2306 2082
rect 2326 2078 2330 2082
rect 2342 2078 2346 2082
rect 2246 1988 2250 1992
rect 2286 2058 2290 2062
rect 2302 2058 2306 2062
rect 2278 2008 2282 2012
rect 2270 1978 2274 1982
rect 2230 1958 2234 1962
rect 2270 1958 2274 1962
rect 2406 2078 2410 2082
rect 2382 2038 2386 2042
rect 2390 2038 2394 2042
rect 2478 2168 2482 2172
rect 2494 2158 2498 2162
rect 2502 2158 2506 2162
rect 2478 2138 2482 2142
rect 2470 2128 2474 2132
rect 2518 2128 2522 2132
rect 2558 2218 2562 2222
rect 2622 2238 2626 2242
rect 2622 2218 2626 2222
rect 2614 2208 2618 2212
rect 2534 2158 2538 2162
rect 2550 2118 2554 2122
rect 2502 2108 2506 2112
rect 2526 2108 2530 2112
rect 2566 2128 2570 2132
rect 2478 2088 2482 2092
rect 2582 2088 2586 2092
rect 2606 2088 2610 2092
rect 2454 2068 2458 2072
rect 2470 2068 2474 2072
rect 2326 2008 2330 2012
rect 2374 2008 2378 2012
rect 2406 2008 2410 2012
rect 2294 1998 2298 2002
rect 2350 1998 2354 2002
rect 2326 1968 2330 1972
rect 2334 1958 2338 1962
rect 2366 1958 2370 1962
rect 2230 1948 2234 1952
rect 2270 1948 2274 1952
rect 2302 1948 2306 1952
rect 2054 1938 2058 1942
rect 2110 1938 2114 1942
rect 2198 1938 2202 1942
rect 2246 1938 2250 1942
rect 2254 1928 2258 1932
rect 2286 1928 2290 1932
rect 2030 1918 2034 1922
rect 2246 1918 2250 1922
rect 2254 1918 2258 1922
rect 1934 1908 1938 1912
rect 1882 1903 1886 1907
rect 1889 1903 1893 1907
rect 1870 1888 1874 1892
rect 1862 1878 1866 1882
rect 1894 1878 1898 1882
rect 1950 1878 1954 1882
rect 1966 1878 1970 1882
rect 1934 1868 1938 1872
rect 1958 1868 1962 1872
rect 1710 1848 1714 1852
rect 1894 1828 1898 1832
rect 1814 1818 1818 1822
rect 1710 1798 1714 1802
rect 1694 1788 1698 1792
rect 1742 1778 1746 1782
rect 1782 1778 1786 1782
rect 1694 1758 1698 1762
rect 1830 1798 1834 1802
rect 1750 1758 1754 1762
rect 1798 1758 1802 1762
rect 1910 1848 1914 1852
rect 1958 1838 1962 1842
rect 1918 1778 1922 1782
rect 1934 1768 1938 1772
rect 1958 1758 1962 1762
rect 1726 1748 1730 1752
rect 1838 1748 1842 1752
rect 1902 1748 1906 1752
rect 1950 1748 1954 1752
rect 1830 1738 1834 1742
rect 1638 1668 1642 1672
rect 1678 1668 1682 1672
rect 1566 1658 1570 1662
rect 1574 1618 1578 1622
rect 1630 1598 1634 1602
rect 1598 1578 1602 1582
rect 1750 1728 1754 1732
rect 1758 1728 1762 1732
rect 1782 1718 1786 1722
rect 1774 1708 1778 1712
rect 1814 1728 1818 1732
rect 1838 1728 1842 1732
rect 1910 1728 1914 1732
rect 1918 1728 1922 1732
rect 1926 1728 1930 1732
rect 1854 1718 1858 1722
rect 1790 1698 1794 1702
rect 1806 1698 1810 1702
rect 1838 1698 1842 1702
rect 1766 1688 1770 1692
rect 1838 1688 1842 1692
rect 1726 1678 1730 1682
rect 1814 1678 1818 1682
rect 1854 1678 1858 1682
rect 1766 1668 1770 1672
rect 1774 1668 1778 1672
rect 1846 1668 1850 1672
rect 1782 1658 1786 1662
rect 1814 1658 1818 1662
rect 1822 1658 1826 1662
rect 1846 1658 1850 1662
rect 1758 1618 1762 1622
rect 1734 1588 1738 1592
rect 1710 1568 1714 1572
rect 1462 1548 1466 1552
rect 1558 1548 1562 1552
rect 1606 1548 1610 1552
rect 1630 1548 1634 1552
rect 1382 1538 1386 1542
rect 1430 1538 1434 1542
rect 1326 1528 1330 1532
rect 1446 1528 1450 1532
rect 1494 1528 1498 1532
rect 1286 1508 1290 1512
rect 1302 1478 1306 1482
rect 1342 1508 1346 1512
rect 1542 1518 1546 1522
rect 1526 1508 1530 1512
rect 1398 1498 1402 1502
rect 1502 1498 1506 1502
rect 1526 1498 1530 1502
rect 1358 1488 1362 1492
rect 1342 1478 1346 1482
rect 1318 1468 1322 1472
rect 1366 1468 1370 1472
rect 1270 1448 1274 1452
rect 1222 1398 1226 1402
rect 1310 1388 1314 1392
rect 1206 1348 1210 1352
rect 1246 1348 1250 1352
rect 1102 1298 1106 1302
rect 1142 1298 1146 1302
rect 1030 1258 1034 1262
rect 998 1248 1002 1252
rect 1022 1198 1026 1202
rect 1126 1288 1130 1292
rect 1142 1288 1146 1292
rect 1110 1268 1114 1272
rect 1150 1278 1154 1282
rect 1158 1268 1162 1272
rect 1182 1268 1186 1272
rect 1262 1318 1266 1322
rect 1254 1298 1258 1302
rect 1086 1258 1090 1262
rect 1134 1258 1138 1262
rect 1110 1228 1114 1232
rect 1054 1158 1058 1162
rect 990 1148 994 1152
rect 1014 1148 1018 1152
rect 1046 1148 1050 1152
rect 1078 1148 1082 1152
rect 990 1138 994 1142
rect 1030 1138 1034 1142
rect 1086 1138 1090 1142
rect 1030 1128 1034 1132
rect 1102 1128 1106 1132
rect 974 1088 978 1092
rect 982 1088 986 1092
rect 974 1078 978 1082
rect 718 1058 722 1062
rect 750 1058 754 1062
rect 774 1058 778 1062
rect 934 1058 938 1062
rect 678 1038 682 1042
rect 630 1028 634 1032
rect 574 998 578 1002
rect 958 1068 962 1072
rect 998 1068 1002 1072
rect 982 1058 986 1062
rect 1022 1098 1026 1102
rect 1086 1098 1090 1102
rect 1014 1068 1018 1072
rect 1030 1078 1034 1082
rect 1030 1058 1034 1062
rect 902 1048 906 1052
rect 966 1048 970 1052
rect 990 1048 994 1052
rect 926 1038 930 1042
rect 950 998 954 1002
rect 998 998 1002 1002
rect 670 948 674 952
rect 702 948 706 952
rect 750 948 754 952
rect 806 948 810 952
rect 910 948 914 952
rect 1030 948 1034 952
rect 550 888 554 892
rect 534 878 538 882
rect 558 878 562 882
rect 398 858 402 862
rect 430 858 434 862
rect 478 858 482 862
rect 406 848 410 852
rect 374 838 378 842
rect 366 818 370 822
rect 390 818 394 822
rect 346 803 350 807
rect 353 803 357 807
rect 374 768 378 772
rect 422 838 426 842
rect 422 768 426 772
rect 342 728 346 732
rect 326 688 330 692
rect 390 728 394 732
rect 494 808 498 812
rect 510 808 514 812
rect 486 748 490 752
rect 454 738 458 742
rect 462 738 466 742
rect 486 738 490 742
rect 502 738 506 742
rect 422 718 426 722
rect 406 708 410 712
rect 406 698 410 702
rect 382 688 386 692
rect 326 678 330 682
rect 358 678 362 682
rect 398 668 402 672
rect 390 658 394 662
rect 346 603 350 607
rect 353 603 357 607
rect 398 648 402 652
rect 422 688 426 692
rect 414 668 418 672
rect 446 678 450 682
rect 310 588 314 592
rect 366 568 370 572
rect 398 568 402 572
rect 278 548 282 552
rect 278 538 282 542
rect 366 538 370 542
rect 390 538 394 542
rect 334 518 338 522
rect 470 728 474 732
rect 462 708 466 712
rect 454 668 458 672
rect 422 658 426 662
rect 422 558 426 562
rect 438 568 442 572
rect 446 568 450 572
rect 430 538 434 542
rect 406 528 410 532
rect 414 528 418 532
rect 366 498 370 502
rect 382 498 386 502
rect 398 498 402 502
rect 422 518 426 522
rect 430 518 434 522
rect 422 508 426 512
rect 302 488 306 492
rect 294 478 298 482
rect 286 468 290 472
rect 230 458 234 462
rect 262 458 266 462
rect 38 358 42 362
rect 86 358 90 362
rect 142 328 146 332
rect 70 298 74 302
rect 86 298 90 302
rect 70 278 74 282
rect 110 208 114 212
rect 174 288 178 292
rect 182 258 186 262
rect 118 188 122 192
rect 158 188 162 192
rect 6 148 10 152
rect 86 148 90 152
rect 38 138 42 142
rect 166 148 170 152
rect 134 108 138 112
rect 118 88 122 92
rect 6 48 10 52
rect 222 218 226 222
rect 198 148 202 152
rect 238 448 242 452
rect 262 448 266 452
rect 262 438 266 442
rect 326 468 330 472
rect 398 468 402 472
rect 414 468 418 472
rect 294 448 298 452
rect 470 668 474 672
rect 486 668 490 672
rect 478 658 482 662
rect 654 918 658 922
rect 574 888 578 892
rect 590 888 594 892
rect 654 868 658 872
rect 1102 1078 1106 1082
rect 1126 1148 1130 1152
rect 1166 1198 1170 1202
rect 1182 1198 1186 1202
rect 1190 1168 1194 1172
rect 1190 1158 1194 1162
rect 1158 1138 1162 1142
rect 1158 1118 1162 1122
rect 1166 1098 1170 1102
rect 1126 1078 1130 1082
rect 1150 1078 1154 1082
rect 1094 1038 1098 1042
rect 1110 1058 1114 1062
rect 1270 1248 1274 1252
rect 1246 1138 1250 1142
rect 1334 1458 1338 1462
rect 1362 1403 1366 1407
rect 1369 1403 1373 1407
rect 1382 1388 1386 1392
rect 1350 1328 1354 1332
rect 1366 1328 1370 1332
rect 1390 1318 1394 1322
rect 1446 1488 1450 1492
rect 1406 1448 1410 1452
rect 1462 1418 1466 1422
rect 1446 1408 1450 1412
rect 1478 1388 1482 1392
rect 1446 1378 1450 1382
rect 1486 1368 1490 1372
rect 1510 1368 1514 1372
rect 1414 1358 1418 1362
rect 1438 1358 1442 1362
rect 1406 1348 1410 1352
rect 1422 1348 1426 1352
rect 1438 1328 1442 1332
rect 1454 1348 1458 1352
rect 1502 1358 1506 1362
rect 1470 1318 1474 1322
rect 1446 1308 1450 1312
rect 1446 1298 1450 1302
rect 1470 1298 1474 1302
rect 1398 1288 1402 1292
rect 1358 1278 1362 1282
rect 1390 1268 1394 1272
rect 1362 1203 1366 1207
rect 1369 1203 1373 1207
rect 1390 1168 1394 1172
rect 1406 1278 1410 1282
rect 1454 1278 1458 1282
rect 1406 1258 1410 1262
rect 1438 1258 1442 1262
rect 1446 1178 1450 1182
rect 1414 1158 1418 1162
rect 1766 1558 1770 1562
rect 1798 1548 1802 1552
rect 1726 1528 1730 1532
rect 1558 1468 1562 1472
rect 1534 1458 1538 1462
rect 1550 1458 1554 1462
rect 1582 1518 1586 1522
rect 1742 1498 1746 1502
rect 1654 1488 1658 1492
rect 1790 1488 1794 1492
rect 1806 1488 1810 1492
rect 1870 1708 1874 1712
rect 1882 1703 1886 1707
rect 1889 1703 1893 1707
rect 1894 1688 1898 1692
rect 1870 1678 1874 1682
rect 1878 1678 1882 1682
rect 1862 1638 1866 1642
rect 1870 1638 1874 1642
rect 1846 1578 1850 1582
rect 1830 1538 1834 1542
rect 1838 1528 1842 1532
rect 1838 1488 1842 1492
rect 1686 1468 1690 1472
rect 1702 1468 1706 1472
rect 1766 1468 1770 1472
rect 1774 1468 1778 1472
rect 1566 1448 1570 1452
rect 1638 1448 1642 1452
rect 1598 1428 1602 1432
rect 1566 1418 1570 1422
rect 1574 1368 1578 1372
rect 1542 1358 1546 1362
rect 1534 1348 1538 1352
rect 1558 1348 1562 1352
rect 1526 1328 1530 1332
rect 1550 1328 1554 1332
rect 1518 1318 1522 1322
rect 1534 1318 1538 1322
rect 1510 1308 1514 1312
rect 1502 1268 1506 1272
rect 1494 1258 1498 1262
rect 1526 1268 1530 1272
rect 1510 1238 1514 1242
rect 1478 1188 1482 1192
rect 1494 1188 1498 1192
rect 1326 1138 1330 1142
rect 1342 1138 1346 1142
rect 1358 1138 1362 1142
rect 1398 1138 1402 1142
rect 1470 1138 1474 1142
rect 1262 1118 1266 1122
rect 1318 1118 1322 1122
rect 1334 1118 1338 1122
rect 1238 1108 1242 1112
rect 1278 1108 1282 1112
rect 1206 1098 1210 1102
rect 1222 1078 1226 1082
rect 1230 1078 1234 1082
rect 1262 1078 1266 1082
rect 1342 1078 1346 1082
rect 1334 1068 1338 1072
rect 1142 1058 1146 1062
rect 1262 1058 1266 1062
rect 1126 1048 1130 1052
rect 1206 1048 1210 1052
rect 1214 1048 1218 1052
rect 1414 1128 1418 1132
rect 1438 1128 1442 1132
rect 1462 1118 1466 1122
rect 1414 1058 1418 1062
rect 1350 1048 1354 1052
rect 1374 1048 1378 1052
rect 1134 1028 1138 1032
rect 1102 958 1106 962
rect 950 938 954 942
rect 1046 938 1050 942
rect 1046 918 1050 922
rect 822 908 826 912
rect 850 903 854 907
rect 857 903 861 907
rect 742 888 746 892
rect 934 888 938 892
rect 1006 888 1010 892
rect 1022 878 1026 882
rect 854 868 858 872
rect 902 868 906 872
rect 670 818 674 822
rect 566 768 570 772
rect 678 756 682 760
rect 558 738 562 742
rect 638 728 642 732
rect 622 718 626 722
rect 606 708 610 712
rect 582 698 586 702
rect 534 668 538 672
rect 526 658 530 662
rect 510 588 514 592
rect 510 568 514 572
rect 502 558 506 562
rect 462 548 466 552
rect 518 548 522 552
rect 582 658 586 662
rect 638 658 642 662
rect 558 648 562 652
rect 542 588 546 592
rect 550 578 554 582
rect 486 538 490 542
rect 526 538 530 542
rect 446 478 450 482
rect 470 478 474 482
rect 494 488 498 492
rect 462 468 466 472
rect 494 468 498 472
rect 510 468 514 472
rect 342 458 346 462
rect 334 448 338 452
rect 438 448 442 452
rect 318 438 322 442
rect 382 438 386 442
rect 398 438 402 442
rect 346 403 350 407
rect 353 403 357 407
rect 558 568 562 572
rect 454 458 458 462
rect 502 458 506 462
rect 542 458 546 462
rect 518 448 522 452
rect 526 448 530 452
rect 510 438 514 442
rect 310 368 314 372
rect 534 348 538 352
rect 494 338 498 342
rect 358 328 362 332
rect 374 328 378 332
rect 286 288 290 292
rect 286 278 290 282
rect 342 258 346 262
rect 630 568 634 572
rect 758 808 762 812
rect 790 808 794 812
rect 1166 1008 1170 1012
rect 1238 998 1242 1002
rect 1206 988 1210 992
rect 1150 958 1154 962
rect 1198 958 1202 962
rect 1166 948 1170 952
rect 1142 938 1146 942
rect 1182 938 1186 942
rect 1190 908 1194 912
rect 1222 908 1226 912
rect 1198 888 1202 892
rect 1222 888 1226 892
rect 1126 868 1130 872
rect 1134 868 1138 872
rect 1150 868 1154 872
rect 1206 868 1210 872
rect 1278 1008 1282 1012
rect 1262 978 1266 982
rect 1362 1003 1366 1007
rect 1369 1003 1373 1007
rect 1494 1118 1498 1122
rect 1478 1108 1482 1112
rect 1526 1248 1530 1252
rect 1638 1418 1642 1422
rect 1614 1398 1618 1402
rect 1598 1328 1602 1332
rect 1566 1298 1570 1302
rect 1566 1278 1570 1282
rect 1630 1358 1634 1362
rect 1646 1378 1650 1382
rect 1662 1358 1666 1362
rect 1726 1458 1730 1462
rect 1758 1458 1762 1462
rect 1790 1458 1794 1462
rect 1806 1458 1810 1462
rect 1718 1388 1722 1392
rect 1710 1378 1714 1382
rect 1638 1348 1642 1352
rect 1702 1348 1706 1352
rect 1622 1328 1626 1332
rect 1638 1328 1642 1332
rect 1606 1268 1610 1272
rect 1582 1258 1586 1262
rect 1558 1248 1562 1252
rect 1534 1238 1538 1242
rect 1518 1218 1522 1222
rect 1518 1178 1522 1182
rect 1542 1168 1546 1172
rect 1518 1158 1522 1162
rect 1574 1158 1578 1162
rect 1542 1148 1546 1152
rect 1574 1148 1578 1152
rect 1526 1128 1530 1132
rect 1542 1118 1546 1122
rect 1574 1118 1578 1122
rect 1598 1248 1602 1252
rect 1686 1318 1690 1322
rect 1742 1378 1746 1382
rect 1798 1448 1802 1452
rect 1814 1448 1818 1452
rect 1798 1418 1802 1422
rect 1766 1378 1770 1382
rect 1774 1368 1778 1372
rect 1750 1358 1754 1362
rect 1766 1358 1770 1362
rect 1758 1348 1762 1352
rect 1782 1348 1786 1352
rect 1926 1708 1930 1712
rect 1942 1708 1946 1712
rect 1918 1688 1922 1692
rect 1934 1698 1938 1702
rect 1950 1678 1954 1682
rect 1886 1658 1890 1662
rect 1918 1658 1922 1662
rect 1886 1608 1890 1612
rect 2102 1908 2106 1912
rect 2038 1888 2042 1892
rect 2094 1878 2098 1882
rect 2022 1868 2026 1872
rect 2078 1868 2082 1872
rect 1982 1838 1986 1842
rect 1990 1818 1994 1822
rect 2174 1878 2178 1882
rect 2014 1848 2018 1852
rect 2070 1848 2074 1852
rect 2102 1848 2106 1852
rect 2054 1838 2058 1842
rect 2006 1798 2010 1802
rect 2086 1798 2090 1802
rect 1998 1788 2002 1792
rect 2030 1768 2034 1772
rect 1974 1758 1978 1762
rect 1998 1748 2002 1752
rect 1966 1728 1970 1732
rect 2062 1758 2066 1762
rect 2134 1828 2138 1832
rect 2126 1788 2130 1792
rect 2110 1778 2114 1782
rect 2086 1748 2090 1752
rect 2118 1758 2122 1762
rect 2150 1808 2154 1812
rect 2022 1738 2026 1742
rect 2070 1738 2074 1742
rect 2102 1738 2106 1742
rect 2134 1738 2138 1742
rect 1982 1728 1986 1732
rect 1974 1708 1978 1712
rect 1982 1688 1986 1692
rect 2022 1728 2026 1732
rect 2054 1728 2058 1732
rect 2054 1698 2058 1702
rect 2030 1688 2034 1692
rect 2022 1678 2026 1682
rect 1990 1668 1994 1672
rect 2006 1668 2010 1672
rect 2038 1668 2042 1672
rect 2230 1848 2234 1852
rect 2222 1808 2226 1812
rect 2190 1758 2194 1762
rect 2230 1758 2234 1762
rect 2246 1758 2250 1762
rect 2158 1738 2162 1742
rect 2150 1728 2154 1732
rect 2134 1718 2138 1722
rect 2094 1708 2098 1712
rect 2102 1708 2106 1712
rect 2142 1698 2146 1702
rect 2110 1688 2114 1692
rect 2078 1678 2082 1682
rect 2126 1678 2130 1682
rect 2062 1668 2066 1672
rect 1958 1658 1962 1662
rect 1990 1638 1994 1642
rect 1958 1598 1962 1602
rect 1918 1538 1922 1542
rect 1862 1528 1866 1532
rect 1882 1503 1886 1507
rect 1889 1503 1893 1507
rect 2118 1648 2122 1652
rect 2110 1638 2114 1642
rect 2094 1588 2098 1592
rect 2214 1728 2218 1732
rect 2198 1698 2202 1702
rect 2294 1898 2298 1902
rect 2262 1888 2266 1892
rect 2278 1878 2282 1882
rect 2294 1878 2298 1882
rect 2310 1938 2314 1942
rect 2326 1938 2330 1942
rect 2350 1938 2354 1942
rect 2318 1928 2322 1932
rect 2310 1898 2314 1902
rect 2366 1908 2370 1912
rect 2358 1878 2362 1882
rect 2294 1868 2298 1872
rect 2302 1858 2306 1862
rect 2310 1848 2314 1852
rect 2326 1838 2330 1842
rect 2366 1858 2370 1862
rect 2350 1838 2354 1842
rect 2386 2003 2390 2007
rect 2393 2003 2397 2007
rect 2398 1988 2402 1992
rect 2406 1958 2410 1962
rect 2446 2058 2450 2062
rect 2430 2038 2434 2042
rect 2470 2038 2474 2042
rect 2446 1998 2450 2002
rect 2430 1968 2434 1972
rect 2526 2078 2530 2082
rect 2550 2078 2554 2082
rect 2574 2068 2578 2072
rect 2582 2068 2586 2072
rect 2598 2068 2602 2072
rect 2638 2178 2642 2182
rect 2542 2058 2546 2062
rect 2566 2058 2570 2062
rect 2590 2058 2594 2062
rect 2486 2048 2490 2052
rect 2510 2048 2514 2052
rect 2510 1978 2514 1982
rect 2438 1958 2442 1962
rect 2446 1958 2450 1962
rect 2414 1948 2418 1952
rect 2422 1948 2426 1952
rect 2422 1938 2426 1942
rect 2446 1938 2450 1942
rect 2470 1938 2474 1942
rect 2478 1938 2482 1942
rect 2422 1918 2426 1922
rect 2470 1888 2474 1892
rect 2422 1878 2426 1882
rect 2446 1878 2450 1882
rect 2430 1868 2434 1872
rect 2470 1868 2474 1872
rect 2390 1848 2394 1852
rect 2374 1818 2378 1822
rect 2386 1803 2390 1807
rect 2393 1803 2397 1807
rect 2334 1798 2338 1802
rect 2286 1728 2290 1732
rect 2366 1728 2370 1732
rect 2230 1688 2234 1692
rect 2310 1678 2314 1682
rect 2334 1668 2338 1672
rect 2302 1658 2306 1662
rect 2190 1598 2194 1602
rect 2158 1578 2162 1582
rect 1982 1548 1986 1552
rect 2038 1548 2042 1552
rect 2094 1548 2098 1552
rect 2102 1548 2106 1552
rect 1966 1538 1970 1542
rect 2022 1518 2026 1522
rect 1942 1488 1946 1492
rect 1854 1468 1858 1472
rect 1870 1458 1874 1462
rect 1902 1458 1906 1462
rect 1838 1428 1842 1432
rect 1822 1418 1826 1422
rect 1838 1418 1842 1422
rect 1814 1358 1818 1362
rect 1830 1348 1834 1352
rect 1846 1348 1850 1352
rect 1734 1338 1738 1342
rect 1734 1328 1738 1332
rect 1846 1338 1850 1342
rect 1726 1308 1730 1312
rect 1750 1308 1754 1312
rect 1694 1298 1698 1302
rect 1718 1298 1722 1302
rect 1822 1318 1826 1322
rect 1646 1288 1650 1292
rect 1742 1288 1746 1292
rect 1806 1288 1810 1292
rect 1702 1268 1706 1272
rect 1782 1268 1786 1272
rect 1734 1258 1738 1262
rect 1750 1248 1754 1252
rect 1734 1238 1738 1242
rect 1758 1238 1762 1242
rect 1638 1228 1642 1232
rect 1718 1228 1722 1232
rect 1646 1218 1650 1222
rect 1638 1168 1642 1172
rect 1622 1158 1626 1162
rect 1606 1148 1610 1152
rect 1622 1148 1626 1152
rect 1654 1198 1658 1202
rect 1686 1198 1690 1202
rect 1662 1178 1666 1182
rect 1590 1118 1594 1122
rect 1614 1128 1618 1132
rect 1630 1128 1634 1132
rect 1606 1118 1610 1122
rect 1630 1118 1634 1122
rect 1462 1078 1466 1082
rect 1446 1068 1450 1072
rect 1494 1078 1498 1082
rect 1558 1078 1562 1082
rect 1622 1078 1626 1082
rect 1470 1058 1474 1062
rect 1478 1058 1482 1062
rect 1502 1058 1506 1062
rect 1470 1048 1474 1052
rect 1494 1048 1498 1052
rect 1590 1068 1594 1072
rect 1638 1068 1642 1072
rect 1742 1218 1746 1222
rect 1814 1248 1818 1252
rect 1766 1188 1770 1192
rect 1806 1188 1810 1192
rect 1742 1178 1746 1182
rect 1734 1168 1738 1172
rect 1718 1148 1722 1152
rect 1670 1128 1674 1132
rect 1678 1088 1682 1092
rect 1710 1088 1714 1092
rect 1670 1078 1674 1082
rect 1582 1058 1586 1062
rect 1622 1058 1626 1062
rect 1694 1058 1698 1062
rect 1718 1058 1722 1062
rect 1526 1048 1530 1052
rect 1534 1048 1538 1052
rect 1510 1038 1514 1042
rect 1574 1038 1578 1042
rect 1430 1008 1434 1012
rect 1398 998 1402 1002
rect 1550 998 1554 1002
rect 1334 948 1338 952
rect 1390 948 1394 952
rect 1294 908 1298 912
rect 1310 908 1314 912
rect 1310 888 1314 892
rect 1294 878 1298 882
rect 1270 868 1274 872
rect 1078 858 1082 862
rect 1086 858 1090 862
rect 1094 858 1098 862
rect 1198 858 1202 862
rect 1230 858 1234 862
rect 1270 858 1274 862
rect 958 828 962 832
rect 910 818 914 822
rect 862 778 866 782
rect 798 768 802 772
rect 838 768 842 772
rect 774 748 778 752
rect 782 748 786 752
rect 734 728 738 732
rect 702 708 706 712
rect 790 708 794 712
rect 718 678 722 682
rect 718 618 722 622
rect 782 558 786 562
rect 590 548 594 552
rect 734 548 738 552
rect 766 548 770 552
rect 646 528 650 532
rect 630 518 634 522
rect 670 488 674 492
rect 758 478 762 482
rect 686 458 690 462
rect 558 438 562 442
rect 598 438 602 442
rect 574 398 578 402
rect 558 388 562 392
rect 590 358 594 362
rect 550 338 554 342
rect 550 318 554 322
rect 502 308 506 312
rect 518 308 522 312
rect 582 308 586 312
rect 462 288 466 292
rect 478 278 482 282
rect 550 278 554 282
rect 574 278 578 282
rect 422 258 426 262
rect 566 258 570 262
rect 334 248 338 252
rect 374 248 378 252
rect 270 208 274 212
rect 326 178 330 182
rect 262 138 266 142
rect 254 128 258 132
rect 278 118 282 122
rect 254 78 258 82
rect 374 218 378 222
rect 494 208 498 212
rect 346 203 350 207
rect 353 203 357 207
rect 350 158 354 162
rect 606 338 610 342
rect 598 278 602 282
rect 598 258 602 262
rect 518 188 522 192
rect 550 188 554 192
rect 510 138 514 142
rect 486 88 490 92
rect 414 78 418 82
rect 502 78 506 82
rect 590 198 594 202
rect 598 148 602 152
rect 614 168 618 172
rect 606 138 610 142
rect 598 98 602 102
rect 638 408 642 412
rect 630 328 634 332
rect 654 398 658 402
rect 822 758 826 762
rect 830 748 834 752
rect 886 748 890 752
rect 822 738 826 742
rect 814 598 818 602
rect 830 708 834 712
rect 850 703 854 707
rect 857 703 861 707
rect 838 698 842 702
rect 838 588 842 592
rect 846 548 850 552
rect 850 503 854 507
rect 857 503 861 507
rect 822 478 826 482
rect 822 468 826 472
rect 838 468 842 472
rect 854 468 858 472
rect 814 458 818 462
rect 822 448 826 452
rect 822 408 826 412
rect 726 388 730 392
rect 750 388 754 392
rect 662 348 666 352
rect 822 348 826 352
rect 734 338 738 342
rect 750 328 754 332
rect 710 308 714 312
rect 670 268 674 272
rect 662 248 666 252
rect 630 228 634 232
rect 662 198 666 202
rect 670 178 674 182
rect 638 158 642 162
rect 758 268 762 272
rect 862 438 866 442
rect 862 368 866 372
rect 1030 758 1034 762
rect 1126 768 1130 772
rect 1182 848 1186 852
rect 1206 848 1210 852
rect 1166 798 1170 802
rect 1158 778 1162 782
rect 1118 748 1122 752
rect 1182 758 1186 762
rect 1174 748 1178 752
rect 1190 748 1194 752
rect 902 738 906 742
rect 1046 738 1050 742
rect 1166 738 1170 742
rect 1150 718 1154 722
rect 958 698 962 702
rect 974 688 978 692
rect 1150 688 1154 692
rect 1134 678 1138 682
rect 1014 658 1018 662
rect 1078 658 1082 662
rect 894 648 898 652
rect 878 608 882 612
rect 974 648 978 652
rect 902 548 906 552
rect 918 518 922 522
rect 910 498 914 502
rect 1062 618 1066 622
rect 1174 608 1178 612
rect 1142 578 1146 582
rect 1054 568 1058 572
rect 1134 558 1138 562
rect 1006 548 1010 552
rect 974 518 978 522
rect 1150 568 1154 572
rect 1158 568 1162 572
rect 1222 748 1226 752
rect 1230 738 1234 742
rect 1222 728 1226 732
rect 1254 788 1258 792
rect 1254 768 1258 772
rect 1270 738 1274 742
rect 1302 848 1306 852
rect 1454 978 1458 982
rect 1558 978 1562 982
rect 1446 948 1450 952
rect 1566 948 1570 952
rect 1398 938 1402 942
rect 1422 938 1426 942
rect 1494 938 1498 942
rect 1558 938 1562 942
rect 1454 918 1458 922
rect 1430 898 1434 902
rect 1414 868 1418 872
rect 1430 828 1434 832
rect 1470 838 1474 842
rect 1326 818 1330 822
rect 1470 808 1474 812
rect 1362 803 1366 807
rect 1369 803 1373 807
rect 1326 798 1330 802
rect 1422 778 1426 782
rect 1318 758 1322 762
rect 1454 768 1458 772
rect 1238 708 1242 712
rect 1294 708 1298 712
rect 1358 708 1362 712
rect 1262 678 1266 682
rect 1278 678 1282 682
rect 1318 678 1322 682
rect 1342 678 1346 682
rect 1238 658 1242 662
rect 1238 648 1242 652
rect 1310 668 1314 672
rect 1342 668 1346 672
rect 1398 688 1402 692
rect 1374 678 1378 682
rect 1406 678 1410 682
rect 1414 668 1418 672
rect 1542 928 1546 932
rect 1526 898 1530 902
rect 1510 868 1514 872
rect 1534 868 1538 872
rect 1494 798 1498 802
rect 1518 858 1522 862
rect 1510 838 1514 842
rect 1510 758 1514 762
rect 1558 878 1562 882
rect 1590 998 1594 1002
rect 1630 1038 1634 1042
rect 1646 1018 1650 1022
rect 1630 1008 1634 1012
rect 1638 1008 1642 1012
rect 1686 998 1690 1002
rect 1646 978 1650 982
rect 1638 968 1642 972
rect 1598 958 1602 962
rect 1598 938 1602 942
rect 1630 928 1634 932
rect 1598 888 1602 892
rect 1590 868 1594 872
rect 1654 958 1658 962
rect 1686 958 1690 962
rect 1774 1158 1778 1162
rect 1750 1148 1754 1152
rect 1782 1138 1786 1142
rect 1798 1128 1802 1132
rect 1726 1048 1730 1052
rect 1694 948 1698 952
rect 1662 928 1666 932
rect 1686 928 1690 932
rect 1662 868 1666 872
rect 1678 878 1682 882
rect 1574 858 1578 862
rect 1598 858 1602 862
rect 1614 858 1618 862
rect 1646 858 1650 862
rect 1670 858 1674 862
rect 1574 848 1578 852
rect 1622 848 1626 852
rect 1630 848 1634 852
rect 1526 838 1530 842
rect 1614 838 1618 842
rect 1614 818 1618 822
rect 1550 758 1554 762
rect 1582 758 1586 762
rect 1598 758 1602 762
rect 1518 748 1522 752
rect 1550 748 1554 752
rect 1574 748 1578 752
rect 1510 738 1514 742
rect 1542 738 1546 742
rect 1502 728 1506 732
rect 1606 728 1610 732
rect 1462 718 1466 722
rect 1286 658 1290 662
rect 1406 658 1410 662
rect 1438 658 1442 662
rect 1310 648 1314 652
rect 1326 648 1330 652
rect 1350 648 1354 652
rect 1262 638 1266 642
rect 1254 608 1258 612
rect 1238 598 1242 602
rect 1206 558 1210 562
rect 1126 548 1130 552
rect 1142 548 1146 552
rect 1182 548 1186 552
rect 1214 548 1218 552
rect 1070 538 1074 542
rect 1118 538 1122 542
rect 1222 538 1226 542
rect 1030 528 1034 532
rect 1038 528 1042 532
rect 1078 528 1082 532
rect 1110 528 1114 532
rect 1158 528 1162 532
rect 1166 528 1170 532
rect 1198 528 1202 532
rect 1230 528 1234 532
rect 1014 508 1018 512
rect 1022 498 1026 502
rect 886 478 890 482
rect 854 348 858 352
rect 846 338 850 342
rect 870 338 874 342
rect 838 328 842 332
rect 850 303 854 307
rect 857 303 861 307
rect 830 288 834 292
rect 846 278 850 282
rect 750 228 754 232
rect 718 168 722 172
rect 638 148 642 152
rect 694 148 698 152
rect 718 148 722 152
rect 630 138 634 142
rect 686 138 690 142
rect 718 138 722 142
rect 622 88 626 92
rect 310 58 314 62
rect 558 58 562 62
rect 582 58 586 62
rect 630 58 634 62
rect 646 58 650 62
rect 238 48 242 52
rect 262 48 266 52
rect 346 3 350 7
rect 353 3 357 7
rect 750 188 754 192
rect 710 98 714 102
rect 734 98 738 102
rect 734 88 738 92
rect 750 78 754 82
rect 806 168 810 172
rect 902 468 906 472
rect 998 488 1002 492
rect 982 478 986 482
rect 918 448 922 452
rect 950 448 954 452
rect 918 388 922 392
rect 926 368 930 372
rect 942 368 946 372
rect 894 358 898 362
rect 902 348 906 352
rect 1014 388 1018 392
rect 966 378 970 382
rect 1022 368 1026 372
rect 902 338 906 342
rect 998 348 1002 352
rect 926 338 930 342
rect 1006 338 1010 342
rect 934 328 938 332
rect 982 328 986 332
rect 918 288 922 292
rect 982 308 986 312
rect 966 298 970 302
rect 998 298 1002 302
rect 950 278 954 282
rect 982 278 986 282
rect 974 268 978 272
rect 950 258 954 262
rect 966 258 970 262
rect 982 248 986 252
rect 974 228 978 232
rect 958 218 962 222
rect 1022 338 1026 342
rect 1102 518 1106 522
rect 1094 478 1098 482
rect 1078 458 1082 462
rect 1150 498 1154 502
rect 1126 478 1130 482
rect 1134 478 1138 482
rect 1142 478 1146 482
rect 1166 518 1170 522
rect 1174 468 1178 472
rect 1286 608 1290 612
rect 1334 628 1338 632
rect 1302 568 1306 572
rect 1310 568 1314 572
rect 1366 638 1370 642
rect 1362 603 1366 607
rect 1369 603 1373 607
rect 1382 588 1386 592
rect 1350 558 1354 562
rect 1294 548 1298 552
rect 1326 548 1330 552
rect 1366 548 1370 552
rect 1262 538 1266 542
rect 1278 508 1282 512
rect 1270 498 1274 502
rect 1174 458 1178 462
rect 1230 458 1234 462
rect 1278 458 1282 462
rect 1094 428 1098 432
rect 1110 398 1114 402
rect 1070 388 1074 392
rect 1086 388 1090 392
rect 1110 388 1114 392
rect 1094 368 1098 372
rect 1150 368 1154 372
rect 1046 348 1050 352
rect 1126 348 1130 352
rect 1150 348 1154 352
rect 1046 338 1050 342
rect 1038 328 1042 332
rect 1046 318 1050 322
rect 1070 308 1074 312
rect 1022 298 1026 302
rect 1014 278 1018 282
rect 1054 288 1058 292
rect 1126 338 1130 342
rect 1102 328 1106 332
rect 1134 328 1138 332
rect 1078 278 1082 282
rect 1094 278 1098 282
rect 1118 278 1122 282
rect 1038 268 1042 272
rect 1110 268 1114 272
rect 1014 258 1018 262
rect 1022 258 1026 262
rect 1046 258 1050 262
rect 990 238 994 242
rect 1030 238 1034 242
rect 998 218 1002 222
rect 1086 258 1090 262
rect 1094 248 1098 252
rect 1070 238 1074 242
rect 1086 218 1090 222
rect 1062 208 1066 212
rect 902 158 906 162
rect 982 178 986 182
rect 1022 178 1026 182
rect 1070 178 1074 182
rect 982 168 986 172
rect 998 168 1002 172
rect 1030 168 1034 172
rect 1046 168 1050 172
rect 1030 158 1034 162
rect 1054 158 1058 162
rect 990 148 994 152
rect 1006 148 1010 152
rect 1054 148 1058 152
rect 1102 168 1106 172
rect 1166 438 1170 442
rect 1190 438 1194 442
rect 1190 378 1194 382
rect 1198 368 1202 372
rect 1286 448 1290 452
rect 1270 438 1274 442
rect 1214 428 1218 432
rect 1246 428 1250 432
rect 1254 428 1258 432
rect 1182 318 1186 322
rect 1190 308 1194 312
rect 1174 268 1178 272
rect 1142 258 1146 262
rect 1166 258 1170 262
rect 1182 258 1186 262
rect 1246 368 1250 372
rect 1246 348 1250 352
rect 1230 328 1234 332
rect 1278 328 1282 332
rect 1214 298 1218 302
rect 1310 538 1314 542
rect 1350 498 1354 502
rect 1342 478 1346 482
rect 1318 458 1322 462
rect 1342 448 1346 452
rect 1390 558 1394 562
rect 1390 528 1394 532
rect 1398 498 1402 502
rect 1390 488 1394 492
rect 1382 458 1386 462
rect 1326 408 1330 412
rect 1302 378 1306 382
rect 1362 403 1366 407
rect 1369 403 1373 407
rect 1542 708 1546 712
rect 1502 698 1506 702
rect 1534 698 1538 702
rect 1478 688 1482 692
rect 1494 688 1498 692
rect 1494 668 1498 672
rect 1518 668 1522 672
rect 1566 688 1570 692
rect 1678 828 1682 832
rect 1662 818 1666 822
rect 1758 1028 1762 1032
rect 1710 1018 1714 1022
rect 1710 1008 1714 1012
rect 1758 998 1762 1002
rect 1774 1088 1778 1092
rect 1790 1068 1794 1072
rect 1782 1058 1786 1062
rect 1782 978 1786 982
rect 1782 968 1786 972
rect 1742 958 1746 962
rect 1766 958 1770 962
rect 1718 948 1722 952
rect 1766 948 1770 952
rect 1846 1308 1850 1312
rect 1838 1298 1842 1302
rect 1886 1448 1890 1452
rect 1910 1438 1914 1442
rect 1878 1388 1882 1392
rect 1934 1458 1938 1462
rect 1918 1378 1922 1382
rect 1862 1328 1866 1332
rect 2094 1468 2098 1472
rect 2038 1448 2042 1452
rect 2054 1448 2058 1452
rect 2070 1398 2074 1402
rect 2006 1368 2010 1372
rect 1926 1318 1930 1322
rect 1902 1308 1906 1312
rect 1882 1303 1886 1307
rect 1889 1303 1893 1307
rect 1854 1278 1858 1282
rect 1934 1278 1938 1282
rect 1918 1268 1922 1272
rect 1982 1268 1986 1272
rect 1854 1248 1858 1252
rect 2006 1318 2010 1322
rect 2038 1318 2042 1322
rect 2150 1508 2154 1512
rect 2198 1568 2202 1572
rect 2286 1608 2290 1612
rect 2502 1928 2506 1932
rect 2590 2048 2594 2052
rect 2622 2048 2626 2052
rect 2558 2038 2562 2042
rect 2526 1978 2530 1982
rect 2542 1968 2546 1972
rect 2622 2018 2626 2022
rect 2598 1978 2602 1982
rect 2590 1948 2594 1952
rect 2526 1938 2530 1942
rect 2558 1938 2562 1942
rect 2606 1938 2610 1942
rect 2518 1908 2522 1912
rect 2694 2448 2698 2452
rect 2718 2428 2722 2432
rect 2686 2378 2690 2382
rect 2678 2358 2682 2362
rect 2702 2358 2706 2362
rect 2750 2458 2754 2462
rect 2734 2428 2738 2432
rect 2726 2398 2730 2402
rect 2758 2368 2762 2372
rect 2734 2358 2738 2362
rect 2702 2338 2706 2342
rect 2750 2338 2754 2342
rect 2718 2318 2722 2322
rect 2806 2508 2810 2512
rect 2790 2488 2794 2492
rect 2822 2528 2826 2532
rect 2814 2488 2818 2492
rect 2814 2478 2818 2482
rect 2822 2458 2826 2462
rect 2854 2638 2858 2642
rect 2886 2668 2890 2672
rect 2878 2658 2882 2662
rect 2906 2703 2910 2707
rect 2913 2703 2917 2707
rect 2902 2668 2906 2672
rect 2926 2668 2930 2672
rect 2862 2628 2866 2632
rect 2966 2948 2970 2952
rect 3150 3248 3154 3252
rect 3182 3248 3186 3252
rect 3126 3238 3130 3242
rect 3158 3238 3162 3242
rect 3182 3238 3186 3242
rect 3198 3238 3202 3242
rect 3126 3208 3130 3212
rect 3158 3178 3162 3182
rect 3142 3158 3146 3162
rect 3150 3158 3154 3162
rect 3166 3158 3170 3162
rect 3174 3158 3178 3162
rect 3094 3098 3098 3102
rect 3118 3098 3122 3102
rect 3078 3088 3082 3092
rect 3102 3088 3106 3092
rect 3086 3078 3090 3082
rect 3110 3068 3114 3072
rect 3070 3058 3074 3062
rect 3094 3058 3098 3062
rect 3054 3038 3058 3042
rect 3062 3008 3066 3012
rect 3046 2998 3050 3002
rect 2990 2858 2994 2862
rect 3014 2848 3018 2852
rect 3102 2908 3106 2912
rect 3054 2868 3058 2872
rect 3086 2858 3090 2862
rect 3038 2848 3042 2852
rect 3070 2848 3074 2852
rect 3174 3148 3178 3152
rect 3134 3128 3138 3132
rect 3150 3128 3154 3132
rect 3158 3128 3162 3132
rect 3134 3108 3138 3112
rect 3166 3088 3170 3092
rect 3126 3058 3130 3062
rect 3126 3048 3130 3052
rect 3142 3058 3146 3062
rect 3150 3008 3154 3012
rect 3150 2988 3154 2992
rect 3134 2978 3138 2982
rect 3126 2958 3130 2962
rect 3110 2868 3114 2872
rect 3158 2968 3162 2972
rect 3230 3248 3234 3252
rect 3230 3238 3234 3242
rect 3238 3238 3242 3242
rect 3206 3218 3210 3222
rect 3206 3158 3210 3162
rect 3190 3138 3194 3142
rect 3182 3058 3186 3062
rect 3182 2998 3186 3002
rect 3214 3118 3218 3122
rect 3214 3108 3218 3112
rect 3302 3408 3306 3412
rect 3326 3388 3330 3392
rect 3294 3368 3298 3372
rect 3302 3368 3306 3372
rect 3318 3368 3322 3372
rect 3310 3348 3314 3352
rect 3294 3338 3298 3342
rect 3318 3318 3322 3322
rect 3278 3268 3282 3272
rect 3302 3268 3306 3272
rect 3286 3258 3290 3262
rect 3294 3248 3298 3252
rect 3366 3378 3370 3382
rect 3350 3368 3354 3372
rect 3462 3558 3466 3562
rect 3502 3558 3506 3562
rect 3662 3558 3666 3562
rect 3454 3548 3458 3552
rect 3462 3548 3466 3552
rect 3470 3548 3474 3552
rect 3534 3548 3538 3552
rect 3566 3548 3570 3552
rect 3606 3548 3610 3552
rect 3446 3538 3450 3542
rect 3382 3518 3386 3522
rect 3382 3458 3386 3462
rect 3390 3458 3394 3462
rect 3342 3358 3346 3362
rect 3374 3358 3378 3362
rect 3334 3348 3338 3352
rect 3478 3538 3482 3542
rect 3510 3528 3514 3532
rect 3478 3518 3482 3522
rect 3518 3488 3522 3492
rect 3462 3478 3466 3482
rect 3518 3478 3522 3482
rect 3438 3468 3442 3472
rect 3478 3468 3482 3472
rect 3430 3458 3434 3462
rect 3438 3458 3442 3462
rect 3502 3448 3506 3452
rect 3494 3438 3498 3442
rect 3462 3428 3466 3432
rect 3414 3418 3418 3422
rect 3366 3348 3370 3352
rect 3382 3348 3386 3352
rect 3334 3298 3338 3302
rect 3350 3328 3354 3332
rect 3342 3288 3346 3292
rect 3342 3278 3346 3282
rect 3350 3268 3354 3272
rect 3382 3328 3386 3332
rect 3382 3318 3386 3322
rect 3454 3408 3458 3412
rect 3410 3403 3414 3407
rect 3417 3403 3421 3407
rect 3550 3538 3554 3542
rect 3662 3538 3666 3542
rect 3646 3528 3650 3532
rect 3566 3508 3570 3512
rect 3542 3498 3546 3502
rect 3598 3518 3602 3522
rect 3590 3498 3594 3502
rect 3582 3488 3586 3492
rect 3606 3478 3610 3482
rect 3582 3468 3586 3472
rect 3526 3458 3530 3462
rect 3550 3458 3554 3462
rect 3566 3458 3570 3462
rect 3622 3458 3626 3462
rect 3590 3448 3594 3452
rect 3526 3438 3530 3442
rect 3558 3438 3562 3442
rect 3518 3428 3522 3432
rect 3542 3428 3546 3432
rect 3550 3418 3554 3422
rect 3574 3408 3578 3412
rect 3502 3398 3506 3402
rect 3430 3388 3434 3392
rect 3478 3388 3482 3392
rect 3486 3388 3490 3392
rect 3422 3358 3426 3362
rect 3486 3348 3490 3352
rect 3406 3338 3410 3342
rect 3454 3338 3458 3342
rect 3438 3318 3442 3322
rect 3398 3308 3402 3312
rect 3398 3278 3402 3282
rect 3358 3258 3362 3262
rect 3366 3258 3370 3262
rect 3398 3258 3402 3262
rect 3406 3258 3410 3262
rect 3422 3258 3426 3262
rect 3326 3248 3330 3252
rect 3390 3248 3394 3252
rect 3438 3248 3442 3252
rect 3310 3218 3314 3222
rect 3374 3218 3378 3222
rect 3270 3208 3274 3212
rect 3262 3198 3266 3202
rect 3262 3178 3266 3182
rect 3254 3128 3258 3132
rect 3230 3098 3234 3102
rect 3198 3078 3202 3082
rect 3206 3068 3210 3072
rect 3238 3068 3242 3072
rect 3238 3058 3242 3062
rect 3230 3048 3234 3052
rect 3238 3038 3242 3042
rect 3190 2968 3194 2972
rect 3230 2968 3234 2972
rect 3238 2958 3242 2962
rect 3230 2948 3234 2952
rect 3174 2928 3178 2932
rect 3262 3118 3266 3122
rect 3254 3088 3258 3092
rect 3278 3178 3282 3182
rect 3366 3198 3370 3202
rect 3350 3178 3354 3182
rect 3318 3158 3322 3162
rect 3334 3158 3338 3162
rect 3286 3148 3290 3152
rect 3326 3148 3330 3152
rect 3302 3128 3306 3132
rect 3254 3068 3258 3072
rect 3262 3058 3266 3062
rect 3294 3068 3298 3072
rect 3358 3138 3362 3142
rect 3410 3203 3414 3207
rect 3417 3203 3421 3207
rect 3382 3158 3386 3162
rect 3398 3158 3402 3162
rect 3430 3158 3434 3162
rect 3494 3328 3498 3332
rect 3462 3318 3466 3322
rect 3478 3288 3482 3292
rect 3606 3418 3610 3422
rect 3598 3388 3602 3392
rect 3582 3368 3586 3372
rect 3598 3368 3602 3372
rect 3510 3358 3514 3362
rect 3558 3358 3562 3362
rect 3518 3348 3522 3352
rect 3526 3348 3530 3352
rect 3550 3348 3554 3352
rect 3462 3278 3466 3282
rect 3486 3258 3490 3262
rect 3526 3328 3530 3332
rect 3534 3298 3538 3302
rect 3518 3278 3522 3282
rect 3510 3258 3514 3262
rect 3542 3288 3546 3292
rect 3550 3268 3554 3272
rect 3550 3258 3554 3262
rect 3526 3248 3530 3252
rect 3542 3248 3546 3252
rect 3502 3238 3506 3242
rect 3550 3238 3554 3242
rect 3438 3148 3442 3152
rect 3470 3148 3474 3152
rect 3590 3358 3594 3362
rect 3646 3498 3650 3502
rect 3710 3528 3714 3532
rect 3734 3528 3738 3532
rect 3742 3528 3746 3532
rect 3694 3488 3698 3492
rect 3670 3468 3674 3472
rect 3678 3448 3682 3452
rect 3702 3448 3706 3452
rect 3630 3438 3634 3442
rect 3662 3438 3666 3442
rect 3670 3438 3674 3442
rect 3654 3428 3658 3432
rect 3630 3398 3634 3402
rect 3614 3378 3618 3382
rect 3630 3368 3634 3372
rect 3622 3358 3626 3362
rect 3606 3348 3610 3352
rect 3702 3428 3706 3432
rect 3694 3398 3698 3402
rect 3670 3378 3674 3382
rect 3686 3348 3690 3352
rect 3686 3338 3690 3342
rect 3638 3328 3642 3332
rect 3662 3328 3666 3332
rect 3670 3328 3674 3332
rect 3678 3308 3682 3312
rect 3646 3298 3650 3302
rect 3662 3298 3666 3302
rect 3614 3288 3618 3292
rect 3606 3268 3610 3272
rect 3574 3258 3578 3262
rect 3638 3288 3642 3292
rect 3614 3258 3618 3262
rect 3638 3268 3642 3272
rect 3646 3258 3650 3262
rect 3582 3238 3586 3242
rect 3590 3238 3594 3242
rect 3550 3178 3554 3182
rect 3542 3168 3546 3172
rect 3566 3168 3570 3172
rect 3502 3158 3506 3162
rect 3550 3158 3554 3162
rect 3502 3148 3506 3152
rect 3390 3138 3394 3142
rect 3406 3138 3410 3142
rect 3446 3138 3450 3142
rect 3478 3138 3482 3142
rect 3486 3138 3490 3142
rect 3342 3128 3346 3132
rect 3398 3128 3402 3132
rect 3374 3098 3378 3102
rect 3350 3088 3354 3092
rect 3334 3058 3338 3062
rect 3366 3058 3370 3062
rect 3270 3018 3274 3022
rect 3382 3038 3386 3042
rect 3398 3038 3402 3042
rect 3438 3128 3442 3132
rect 3534 3138 3538 3142
rect 3518 3128 3522 3132
rect 3430 3078 3434 3082
rect 3510 3078 3514 3082
rect 3526 3088 3530 3092
rect 3470 3058 3474 3062
rect 3478 3058 3482 3062
rect 3494 3058 3498 3062
rect 3518 3058 3522 3062
rect 3430 3048 3434 3052
rect 3326 3018 3330 3022
rect 3406 3018 3410 3022
rect 3414 3018 3418 3022
rect 3294 3008 3298 3012
rect 3310 3008 3314 3012
rect 3410 3003 3414 3007
rect 3417 3003 3421 3007
rect 3334 2988 3338 2992
rect 3342 2978 3346 2982
rect 3414 2978 3418 2982
rect 3254 2968 3258 2972
rect 3270 2968 3274 2972
rect 3318 2968 3322 2972
rect 3350 2968 3354 2972
rect 3286 2958 3290 2962
rect 3302 2948 3306 2952
rect 3318 2948 3322 2952
rect 3326 2948 3330 2952
rect 3342 2948 3346 2952
rect 3270 2938 3274 2942
rect 3262 2928 3266 2932
rect 3150 2918 3154 2922
rect 3118 2858 3122 2862
rect 3214 2898 3218 2902
rect 3166 2888 3170 2892
rect 3246 2888 3250 2892
rect 3150 2878 3154 2882
rect 3206 2878 3210 2882
rect 3374 2948 3378 2952
rect 3390 2948 3394 2952
rect 3286 2928 3290 2932
rect 3310 2918 3314 2922
rect 3262 2888 3266 2892
rect 3254 2868 3258 2872
rect 3198 2858 3202 2862
rect 3102 2848 3106 2852
rect 3150 2848 3154 2852
rect 2990 2838 2994 2842
rect 3030 2838 3034 2842
rect 3062 2838 3066 2842
rect 3094 2838 3098 2842
rect 3038 2828 3042 2832
rect 3070 2828 3074 2832
rect 3230 2828 3234 2832
rect 2998 2788 3002 2792
rect 3022 2748 3026 2752
rect 3006 2738 3010 2742
rect 2958 2708 2962 2712
rect 3078 2768 3082 2772
rect 3078 2748 3082 2752
rect 3086 2748 3090 2752
rect 3054 2698 3058 2702
rect 3046 2688 3050 2692
rect 2942 2668 2946 2672
rect 3030 2658 3034 2662
rect 2966 2648 2970 2652
rect 3126 2798 3130 2802
rect 3158 2798 3162 2802
rect 3102 2748 3106 2752
rect 3374 2918 3378 2922
rect 3382 2918 3386 2922
rect 3390 2918 3394 2922
rect 3358 2888 3362 2892
rect 3310 2878 3314 2882
rect 3366 2878 3370 2882
rect 3278 2868 3282 2872
rect 3262 2858 3266 2862
rect 3302 2848 3306 2852
rect 3334 2868 3338 2872
rect 3334 2848 3338 2852
rect 3342 2848 3346 2852
rect 3302 2828 3306 2832
rect 3318 2828 3322 2832
rect 3358 2828 3362 2832
rect 3238 2788 3242 2792
rect 3174 2718 3178 2722
rect 3142 2698 3146 2702
rect 3166 2698 3170 2702
rect 3294 2768 3298 2772
rect 3270 2758 3274 2762
rect 3278 2748 3282 2752
rect 3262 2738 3266 2742
rect 3366 2818 3370 2822
rect 3350 2768 3354 2772
rect 3358 2758 3362 2762
rect 3382 2858 3386 2862
rect 3422 2938 3426 2942
rect 3422 2868 3426 2872
rect 3398 2828 3402 2832
rect 3406 2828 3410 2832
rect 3382 2768 3386 2772
rect 3374 2748 3378 2752
rect 3410 2803 3414 2807
rect 3417 2803 3421 2807
rect 3430 2798 3434 2802
rect 3454 3048 3458 3052
rect 3462 3038 3466 3042
rect 3454 3018 3458 3022
rect 3446 2988 3450 2992
rect 3518 3048 3522 3052
rect 3526 3048 3530 3052
rect 3566 3148 3570 3152
rect 3574 3148 3578 3152
rect 3598 3158 3602 3162
rect 3630 3158 3634 3162
rect 3686 3278 3690 3282
rect 3694 3278 3698 3282
rect 3758 3498 3762 3502
rect 3742 3478 3746 3482
rect 3726 3468 3730 3472
rect 3718 3378 3722 3382
rect 3734 3398 3738 3402
rect 3726 3368 3730 3372
rect 3718 3358 3722 3362
rect 3710 3338 3714 3342
rect 3718 3328 3722 3332
rect 3774 3438 3778 3442
rect 3750 3408 3754 3412
rect 3750 3338 3754 3342
rect 3742 3328 3746 3332
rect 3758 3328 3762 3332
rect 3734 3308 3738 3312
rect 3726 3298 3730 3302
rect 3774 3368 3778 3372
rect 3742 3278 3746 3282
rect 3766 3278 3770 3282
rect 3718 3258 3722 3262
rect 3766 3258 3770 3262
rect 3710 3248 3714 3252
rect 3726 3248 3730 3252
rect 3718 3238 3722 3242
rect 3766 3228 3770 3232
rect 3702 3218 3706 3222
rect 3718 3218 3722 3222
rect 3678 3188 3682 3192
rect 3702 3178 3706 3182
rect 3686 3168 3690 3172
rect 3614 3148 3618 3152
rect 3662 3148 3666 3152
rect 3606 3138 3610 3142
rect 3590 3128 3594 3132
rect 3566 3048 3570 3052
rect 3582 3048 3586 3052
rect 3518 3028 3522 3032
rect 3510 3018 3514 3022
rect 3478 2998 3482 3002
rect 3526 3018 3530 3022
rect 3462 2978 3466 2982
rect 3518 2978 3522 2982
rect 3502 2968 3506 2972
rect 3470 2948 3474 2952
rect 3534 2958 3538 2962
rect 3590 3038 3594 3042
rect 3566 2998 3570 3002
rect 3542 2948 3546 2952
rect 3454 2928 3458 2932
rect 3462 2928 3466 2932
rect 3526 2928 3530 2932
rect 3526 2898 3530 2902
rect 3470 2888 3474 2892
rect 3518 2878 3522 2882
rect 3710 3168 3714 3172
rect 3726 3158 3730 3162
rect 3654 3138 3658 3142
rect 3742 3138 3746 3142
rect 3654 3128 3658 3132
rect 3630 3078 3634 3082
rect 3678 3118 3682 3122
rect 3726 3118 3730 3122
rect 3654 3078 3658 3082
rect 3702 3088 3706 3092
rect 3718 3088 3722 3092
rect 3678 3078 3682 3082
rect 3702 3078 3706 3082
rect 3662 3068 3666 3072
rect 3750 3098 3754 3102
rect 3742 3068 3746 3072
rect 3630 3058 3634 3062
rect 3742 3058 3746 3062
rect 3614 2988 3618 2992
rect 3590 2978 3594 2982
rect 3582 2968 3586 2972
rect 3574 2928 3578 2932
rect 3566 2918 3570 2922
rect 3558 2898 3562 2902
rect 3574 2878 3578 2882
rect 3622 2958 3626 2962
rect 3662 3048 3666 3052
rect 3694 3048 3698 3052
rect 3734 3048 3738 3052
rect 3702 3038 3706 3042
rect 3686 3008 3690 3012
rect 3606 2948 3610 2952
rect 3654 2948 3658 2952
rect 3670 2948 3674 2952
rect 3622 2938 3626 2942
rect 3646 2938 3650 2942
rect 3654 2938 3658 2942
rect 3662 2938 3666 2942
rect 3574 2868 3578 2872
rect 3454 2848 3458 2852
rect 3438 2788 3442 2792
rect 3438 2768 3442 2772
rect 3590 2848 3594 2852
rect 3646 2918 3650 2922
rect 3606 2878 3610 2882
rect 3630 2868 3634 2872
rect 3758 2948 3762 2952
rect 3766 2948 3770 2952
rect 3694 2928 3698 2932
rect 3702 2928 3706 2932
rect 3662 2908 3666 2912
rect 3670 2888 3674 2892
rect 3662 2878 3666 2882
rect 3614 2858 3618 2862
rect 3550 2828 3554 2832
rect 3630 2828 3634 2832
rect 3494 2818 3498 2822
rect 3542 2818 3546 2822
rect 3494 2798 3498 2802
rect 3454 2758 3458 2762
rect 3534 2768 3538 2772
rect 3566 2778 3570 2782
rect 3598 2778 3602 2782
rect 3502 2758 3506 2762
rect 3518 2758 3522 2762
rect 3542 2758 3546 2762
rect 3742 2938 3746 2942
rect 3758 2938 3762 2942
rect 3734 2928 3738 2932
rect 3734 2878 3738 2882
rect 3750 2918 3754 2922
rect 3766 2888 3770 2892
rect 3758 2878 3762 2882
rect 3686 2858 3690 2862
rect 3726 2778 3730 2782
rect 3774 2808 3778 2812
rect 3718 2768 3722 2772
rect 3750 2768 3754 2772
rect 3654 2758 3658 2762
rect 3662 2758 3666 2762
rect 3686 2758 3690 2762
rect 3550 2748 3554 2752
rect 3590 2748 3594 2752
rect 3622 2748 3626 2752
rect 3422 2738 3426 2742
rect 3470 2738 3474 2742
rect 3358 2728 3362 2732
rect 3414 2728 3418 2732
rect 3326 2718 3330 2722
rect 3406 2718 3410 2722
rect 3262 2708 3266 2712
rect 3294 2708 3298 2712
rect 3262 2688 3266 2692
rect 3166 2678 3170 2682
rect 3182 2678 3186 2682
rect 3334 2708 3338 2712
rect 3350 2698 3354 2702
rect 3486 2698 3490 2702
rect 3486 2688 3490 2692
rect 3294 2678 3298 2682
rect 3158 2668 3162 2672
rect 3198 2668 3202 2672
rect 3214 2668 3218 2672
rect 3222 2668 3226 2672
rect 3278 2668 3282 2672
rect 3286 2668 3290 2672
rect 3326 2668 3330 2672
rect 3190 2658 3194 2662
rect 3094 2648 3098 2652
rect 3118 2638 3122 2642
rect 3198 2648 3202 2652
rect 3190 2628 3194 2632
rect 3094 2618 3098 2622
rect 2998 2608 3002 2612
rect 2990 2598 2994 2602
rect 2854 2588 2858 2592
rect 2942 2588 2946 2592
rect 2958 2578 2962 2582
rect 2862 2568 2866 2572
rect 2846 2558 2850 2562
rect 2974 2558 2978 2562
rect 2982 2548 2986 2552
rect 2854 2528 2858 2532
rect 3046 2578 3050 2582
rect 3086 2578 3090 2582
rect 3038 2558 3042 2562
rect 3030 2548 3034 2552
rect 2886 2538 2890 2542
rect 2902 2538 2906 2542
rect 2886 2528 2890 2532
rect 2886 2508 2890 2512
rect 2906 2503 2910 2507
rect 2913 2503 2917 2507
rect 2894 2498 2898 2502
rect 2942 2528 2946 2532
rect 3070 2568 3074 2572
rect 3062 2548 3066 2552
rect 3110 2578 3114 2582
rect 3206 2588 3210 2592
rect 3174 2558 3178 2562
rect 3182 2558 3186 2562
rect 3166 2548 3170 2552
rect 3094 2538 3098 2542
rect 3014 2528 3018 2532
rect 3070 2528 3074 2532
rect 3102 2528 3106 2532
rect 2870 2488 2874 2492
rect 2894 2488 2898 2492
rect 2838 2468 2842 2472
rect 2878 2468 2882 2472
rect 2958 2478 2962 2482
rect 2990 2478 2994 2482
rect 3094 2518 3098 2522
rect 3022 2478 3026 2482
rect 2926 2468 2930 2472
rect 2982 2468 2986 2472
rect 3006 2468 3010 2472
rect 2846 2458 2850 2462
rect 2862 2458 2866 2462
rect 2902 2458 2906 2462
rect 2830 2448 2834 2452
rect 2798 2438 2802 2442
rect 2782 2428 2786 2432
rect 2774 2388 2778 2392
rect 2814 2398 2818 2402
rect 2830 2388 2834 2392
rect 2838 2388 2842 2392
rect 2798 2338 2802 2342
rect 2766 2328 2770 2332
rect 2806 2328 2810 2332
rect 2774 2318 2778 2322
rect 2734 2288 2738 2292
rect 2878 2448 2882 2452
rect 2870 2388 2874 2392
rect 2894 2368 2898 2372
rect 2838 2348 2842 2352
rect 2846 2348 2850 2352
rect 2862 2348 2866 2352
rect 2878 2348 2882 2352
rect 2830 2298 2834 2302
rect 2734 2268 2738 2272
rect 2774 2268 2778 2272
rect 2822 2268 2826 2272
rect 2718 2258 2722 2262
rect 2782 2258 2786 2262
rect 2814 2248 2818 2252
rect 2774 2188 2778 2192
rect 2806 2188 2810 2192
rect 2758 2178 2762 2182
rect 2662 2158 2666 2162
rect 2678 2158 2682 2162
rect 2694 2158 2698 2162
rect 2678 2148 2682 2152
rect 2742 2148 2746 2152
rect 2718 2138 2722 2142
rect 2686 2118 2690 2122
rect 2670 2108 2674 2112
rect 2670 2098 2674 2102
rect 2662 2088 2666 2092
rect 2654 2078 2658 2082
rect 2662 2068 2666 2072
rect 2726 2128 2730 2132
rect 2734 2108 2738 2112
rect 2694 2098 2698 2102
rect 2734 2098 2738 2102
rect 2726 2078 2730 2082
rect 2854 2338 2858 2342
rect 2878 2338 2882 2342
rect 2862 2298 2866 2302
rect 2906 2303 2910 2307
rect 2913 2303 2917 2307
rect 2958 2458 2962 2462
rect 2974 2458 2978 2462
rect 2998 2458 3002 2462
rect 2990 2448 2994 2452
rect 3062 2478 3066 2482
rect 3070 2478 3074 2482
rect 3086 2478 3090 2482
rect 3030 2368 3034 2372
rect 2998 2358 3002 2362
rect 2998 2348 3002 2352
rect 3062 2428 3066 2432
rect 3070 2418 3074 2422
rect 3062 2358 3066 2362
rect 2982 2338 2986 2342
rect 3030 2338 3034 2342
rect 3038 2318 3042 2322
rect 3006 2308 3010 2312
rect 2942 2288 2946 2292
rect 2958 2288 2962 2292
rect 2974 2288 2978 2292
rect 2942 2278 2946 2282
rect 3046 2288 3050 2292
rect 3030 2278 3034 2282
rect 3038 2278 3042 2282
rect 3078 2368 3082 2372
rect 3150 2528 3154 2532
rect 3118 2518 3122 2522
rect 3134 2518 3138 2522
rect 3142 2508 3146 2512
rect 3174 2498 3178 2502
rect 3118 2488 3122 2492
rect 3110 2468 3114 2472
rect 3150 2478 3154 2482
rect 3142 2468 3146 2472
rect 3078 2358 3082 2362
rect 3086 2358 3090 2362
rect 3198 2478 3202 2482
rect 3230 2648 3234 2652
rect 3230 2618 3234 2622
rect 3214 2578 3218 2582
rect 3254 2608 3258 2612
rect 3254 2578 3258 2582
rect 3222 2558 3226 2562
rect 3238 2558 3242 2562
rect 3262 2558 3266 2562
rect 3334 2648 3338 2652
rect 3342 2648 3346 2652
rect 3318 2568 3322 2572
rect 3326 2568 3330 2572
rect 3326 2548 3330 2552
rect 3222 2538 3226 2542
rect 3222 2518 3226 2522
rect 3230 2488 3234 2492
rect 3246 2488 3250 2492
rect 3246 2468 3250 2472
rect 3134 2438 3138 2442
rect 3166 2438 3170 2442
rect 3182 2438 3186 2442
rect 3102 2418 3106 2422
rect 3126 2418 3130 2422
rect 3118 2358 3122 2362
rect 3166 2418 3170 2422
rect 3262 2518 3266 2522
rect 3342 2558 3346 2562
rect 3350 2558 3354 2562
rect 3382 2648 3386 2652
rect 3374 2608 3378 2612
rect 3366 2538 3370 2542
rect 3310 2508 3314 2512
rect 3262 2488 3266 2492
rect 3302 2488 3306 2492
rect 3270 2478 3274 2482
rect 3214 2438 3218 2442
rect 3262 2388 3266 2392
rect 3206 2378 3210 2382
rect 3230 2368 3234 2372
rect 3158 2358 3162 2362
rect 3166 2348 3170 2352
rect 3214 2348 3218 2352
rect 3118 2338 3122 2342
rect 3166 2338 3170 2342
rect 3190 2338 3194 2342
rect 3246 2338 3250 2342
rect 3078 2318 3082 2322
rect 3070 2298 3074 2302
rect 2886 2268 2890 2272
rect 2950 2268 2954 2272
rect 2998 2268 3002 2272
rect 3022 2268 3026 2272
rect 3046 2268 3050 2272
rect 2878 2258 2882 2262
rect 2838 2178 2842 2182
rect 2814 2168 2818 2172
rect 2822 2148 2826 2152
rect 2790 2138 2794 2142
rect 2846 2138 2850 2142
rect 2782 2128 2786 2132
rect 2822 2128 2826 2132
rect 2766 2118 2770 2122
rect 2862 2188 2866 2192
rect 2862 2148 2866 2152
rect 2854 2098 2858 2102
rect 2822 2088 2826 2092
rect 2806 2078 2810 2082
rect 2758 2068 2762 2072
rect 2702 2058 2706 2062
rect 2662 2048 2666 2052
rect 2662 2038 2666 2042
rect 2670 2038 2674 2042
rect 2694 2038 2698 2042
rect 2638 1968 2642 1972
rect 2958 2258 2962 2262
rect 2990 2258 2994 2262
rect 2934 2248 2938 2252
rect 2982 2248 2986 2252
rect 2998 2248 3002 2252
rect 2910 2208 2914 2212
rect 2902 2188 2906 2192
rect 3022 2188 3026 2192
rect 2902 2148 2906 2152
rect 2950 2138 2954 2142
rect 3182 2328 3186 2332
rect 3158 2318 3162 2322
rect 3134 2308 3138 2312
rect 3110 2278 3114 2282
rect 3046 2258 3050 2262
rect 3102 2258 3106 2262
rect 3118 2258 3122 2262
rect 3102 2238 3106 2242
rect 3070 2218 3074 2222
rect 3102 2198 3106 2202
rect 3126 2248 3130 2252
rect 3134 2248 3138 2252
rect 3166 2248 3170 2252
rect 3126 2168 3130 2172
rect 3110 2158 3114 2162
rect 3126 2158 3130 2162
rect 3038 2138 3042 2142
rect 3046 2138 3050 2142
rect 3078 2138 3082 2142
rect 3110 2138 3114 2142
rect 2886 2128 2890 2132
rect 2966 2128 2970 2132
rect 3030 2128 3034 2132
rect 3022 2108 3026 2112
rect 2906 2103 2910 2107
rect 2913 2103 2917 2107
rect 2990 2098 2994 2102
rect 2966 2088 2970 2092
rect 2950 2078 2954 2082
rect 2942 2058 2946 2062
rect 2958 2058 2962 2062
rect 2934 2048 2938 2052
rect 2894 2028 2898 2032
rect 2742 2018 2746 2022
rect 2806 2018 2810 2022
rect 2830 2018 2834 2022
rect 2718 1998 2722 2002
rect 2742 1998 2746 2002
rect 2718 1968 2722 1972
rect 2654 1938 2658 1942
rect 2686 1928 2690 1932
rect 2718 1948 2722 1952
rect 2702 1938 2706 1942
rect 2710 1938 2714 1942
rect 2574 1918 2578 1922
rect 2694 1918 2698 1922
rect 2534 1908 2538 1912
rect 2526 1898 2530 1902
rect 2502 1868 2506 1872
rect 2734 1918 2738 1922
rect 2726 1898 2730 1902
rect 2550 1868 2554 1872
rect 2662 1868 2666 1872
rect 2494 1858 2498 1862
rect 2518 1858 2522 1862
rect 2414 1848 2418 1852
rect 2454 1848 2458 1852
rect 2526 1848 2530 1852
rect 2486 1818 2490 1822
rect 2462 1758 2466 1762
rect 2510 1758 2514 1762
rect 2406 1708 2410 1712
rect 2366 1688 2370 1692
rect 2366 1678 2370 1682
rect 2486 1738 2490 1742
rect 2518 1738 2522 1742
rect 2478 1728 2482 1732
rect 2470 1698 2474 1702
rect 2470 1688 2474 1692
rect 2414 1658 2418 1662
rect 2358 1618 2362 1622
rect 2386 1603 2390 1607
rect 2393 1603 2397 1607
rect 2350 1558 2354 1562
rect 2438 1558 2442 1562
rect 2454 1558 2458 1562
rect 2214 1548 2218 1552
rect 2246 1528 2250 1532
rect 2278 1528 2282 1532
rect 2294 1528 2298 1532
rect 2246 1498 2250 1502
rect 2078 1348 2082 1352
rect 2070 1298 2074 1302
rect 2046 1268 2050 1272
rect 2126 1438 2130 1442
rect 2134 1368 2138 1372
rect 2118 1358 2122 1362
rect 2134 1348 2138 1352
rect 2126 1328 2130 1332
rect 2230 1458 2234 1462
rect 2246 1458 2250 1462
rect 2190 1398 2194 1402
rect 2214 1398 2218 1402
rect 2230 1398 2234 1402
rect 2190 1368 2194 1372
rect 2158 1358 2162 1362
rect 2166 1338 2170 1342
rect 2198 1338 2202 1342
rect 2182 1328 2186 1332
rect 2206 1328 2210 1332
rect 2182 1308 2186 1312
rect 2014 1258 2018 1262
rect 2046 1258 2050 1262
rect 2086 1258 2090 1262
rect 2102 1258 2106 1262
rect 1990 1238 1994 1242
rect 2006 1228 2010 1232
rect 2022 1218 2026 1222
rect 1902 1208 1906 1212
rect 1934 1188 1938 1192
rect 1926 1178 1930 1182
rect 1918 1158 1922 1162
rect 1862 1148 1866 1152
rect 1822 1138 1826 1142
rect 1862 1128 1866 1132
rect 1902 1118 1906 1122
rect 2054 1198 2058 1202
rect 2142 1168 2146 1172
rect 2038 1148 2042 1152
rect 2070 1138 2074 1142
rect 2022 1128 2026 1132
rect 2038 1118 2042 1122
rect 1870 1108 1874 1112
rect 1926 1108 1930 1112
rect 1882 1103 1886 1107
rect 1889 1103 1893 1107
rect 1998 1108 2002 1112
rect 2038 1108 2042 1112
rect 1830 1098 1834 1102
rect 1942 1098 1946 1102
rect 1894 1088 1898 1092
rect 1998 1088 2002 1092
rect 1878 1078 1882 1082
rect 1998 1068 2002 1072
rect 2022 1058 2026 1062
rect 2110 1118 2114 1122
rect 2166 1238 2170 1242
rect 2150 1158 2154 1162
rect 2238 1388 2242 1392
rect 2310 1468 2314 1472
rect 2542 1838 2546 1842
rect 2614 1858 2618 1862
rect 2606 1848 2610 1852
rect 2574 1818 2578 1822
rect 2550 1798 2554 1802
rect 2542 1748 2546 1752
rect 2550 1748 2554 1752
rect 2582 1768 2586 1772
rect 2678 1798 2682 1802
rect 2646 1768 2650 1772
rect 2638 1758 2642 1762
rect 2574 1748 2578 1752
rect 2622 1748 2626 1752
rect 2550 1738 2554 1742
rect 2558 1738 2562 1742
rect 2582 1738 2586 1742
rect 2542 1688 2546 1692
rect 2574 1728 2578 1732
rect 2550 1678 2554 1682
rect 2598 1698 2602 1702
rect 2590 1678 2594 1682
rect 2574 1668 2578 1672
rect 2582 1658 2586 1662
rect 2566 1648 2570 1652
rect 2542 1618 2546 1622
rect 2518 1608 2522 1612
rect 2454 1548 2458 1552
rect 2510 1548 2514 1552
rect 2590 1558 2594 1562
rect 2702 1768 2706 1772
rect 2718 1768 2722 1772
rect 2878 2008 2882 2012
rect 2862 1988 2866 1992
rect 2790 1968 2794 1972
rect 2814 1958 2818 1962
rect 2862 1958 2866 1962
rect 2766 1948 2770 1952
rect 2758 1938 2762 1942
rect 2766 1928 2770 1932
rect 2782 1918 2786 1922
rect 2782 1898 2786 1902
rect 2894 1958 2898 1962
rect 2862 1948 2866 1952
rect 2886 1948 2890 1952
rect 2926 1948 2930 1952
rect 2798 1938 2802 1942
rect 2854 1938 2858 1942
rect 2950 1958 2954 1962
rect 2950 1948 2954 1952
rect 2958 1938 2962 1942
rect 2806 1928 2810 1932
rect 2838 1918 2842 1922
rect 2814 1908 2818 1912
rect 2790 1888 2794 1892
rect 2790 1868 2794 1872
rect 2750 1848 2754 1852
rect 2662 1758 2666 1762
rect 2726 1758 2730 1762
rect 2678 1748 2682 1752
rect 2742 1748 2746 1752
rect 2670 1738 2674 1742
rect 2694 1738 2698 1742
rect 2710 1738 2714 1742
rect 2726 1738 2730 1742
rect 2638 1728 2642 1732
rect 2606 1618 2610 1622
rect 2654 1698 2658 1702
rect 2646 1678 2650 1682
rect 2670 1708 2674 1712
rect 2686 1708 2690 1712
rect 2678 1688 2682 1692
rect 2638 1668 2642 1672
rect 2662 1668 2666 1672
rect 2630 1658 2634 1662
rect 2646 1658 2650 1662
rect 2702 1698 2706 1702
rect 2710 1698 2714 1702
rect 2726 1678 2730 1682
rect 2670 1648 2674 1652
rect 2662 1638 2666 1642
rect 2646 1588 2650 1592
rect 2622 1568 2626 1572
rect 2550 1538 2554 1542
rect 2574 1538 2578 1542
rect 2598 1538 2602 1542
rect 2454 1528 2458 1532
rect 2526 1528 2530 1532
rect 2350 1508 2354 1512
rect 2366 1498 2370 1502
rect 2390 1498 2394 1502
rect 2334 1468 2338 1472
rect 2366 1468 2370 1472
rect 2446 1468 2450 1472
rect 2326 1458 2330 1462
rect 2302 1448 2306 1452
rect 2254 1398 2258 1402
rect 2318 1398 2322 1402
rect 2294 1368 2298 1372
rect 2398 1458 2402 1462
rect 2358 1438 2362 1442
rect 2430 1418 2434 1422
rect 2358 1408 2362 1412
rect 2386 1403 2390 1407
rect 2393 1403 2397 1407
rect 2358 1388 2362 1392
rect 2382 1368 2386 1372
rect 2414 1368 2418 1372
rect 2270 1358 2274 1362
rect 2286 1358 2290 1362
rect 2246 1328 2250 1332
rect 2230 1268 2234 1272
rect 2350 1348 2354 1352
rect 2286 1338 2290 1342
rect 2326 1338 2330 1342
rect 2358 1338 2362 1342
rect 2326 1328 2330 1332
rect 2254 1318 2258 1322
rect 2318 1318 2322 1322
rect 2302 1298 2306 1302
rect 2262 1288 2266 1292
rect 2286 1288 2290 1292
rect 2294 1288 2298 1292
rect 2246 1268 2250 1272
rect 2222 1218 2226 1222
rect 2238 1208 2242 1212
rect 2270 1258 2274 1262
rect 2334 1298 2338 1302
rect 2406 1328 2410 1332
rect 2398 1318 2402 1322
rect 2374 1308 2378 1312
rect 2398 1308 2402 1312
rect 2374 1288 2378 1292
rect 2398 1278 2402 1282
rect 2358 1268 2362 1272
rect 2382 1268 2386 1272
rect 2302 1238 2306 1242
rect 2310 1238 2314 1242
rect 2294 1208 2298 1212
rect 2254 1178 2258 1182
rect 2214 1128 2218 1132
rect 2246 1128 2250 1132
rect 2158 1118 2162 1122
rect 2214 1118 2218 1122
rect 2086 1088 2090 1092
rect 2110 1088 2114 1092
rect 2054 1078 2058 1082
rect 2094 1078 2098 1082
rect 2070 1068 2074 1072
rect 2086 1058 2090 1062
rect 1822 1028 1826 1032
rect 1894 1048 1898 1052
rect 2022 1048 2026 1052
rect 2078 1048 2082 1052
rect 1854 998 1858 1002
rect 1806 948 1810 952
rect 1830 948 1834 952
rect 1886 948 1890 952
rect 2030 1038 2034 1042
rect 2102 1038 2106 1042
rect 2062 1018 2066 1022
rect 1974 998 1978 1002
rect 1982 998 1986 1002
rect 1910 968 1914 972
rect 1958 958 1962 962
rect 2198 1078 2202 1082
rect 2126 1038 2130 1042
rect 2150 1058 2154 1062
rect 2134 1018 2138 1022
rect 2150 1018 2154 1022
rect 2174 1068 2178 1072
rect 2190 1068 2194 1072
rect 2182 1058 2186 1062
rect 2158 998 2162 1002
rect 2166 978 2170 982
rect 2118 958 2122 962
rect 2150 958 2154 962
rect 1926 948 1930 952
rect 1950 948 1954 952
rect 1982 948 1986 952
rect 2054 948 2058 952
rect 1758 938 1762 942
rect 1806 938 1810 942
rect 1838 938 1842 942
rect 1854 938 1858 942
rect 1862 938 1866 942
rect 1950 938 1954 942
rect 1974 938 1978 942
rect 1702 928 1706 932
rect 1734 928 1738 932
rect 1694 858 1698 862
rect 1686 768 1690 772
rect 1638 748 1642 752
rect 1678 748 1682 752
rect 1670 738 1674 742
rect 1630 728 1634 732
rect 1670 698 1674 702
rect 1686 698 1690 702
rect 1574 678 1578 682
rect 1622 678 1626 682
rect 1566 668 1570 672
rect 1510 648 1514 652
rect 1438 598 1442 602
rect 1430 558 1434 562
rect 1502 598 1506 602
rect 1486 588 1490 592
rect 1486 578 1490 582
rect 1606 668 1610 672
rect 1614 658 1618 662
rect 1614 628 1618 632
rect 1590 618 1594 622
rect 1574 608 1578 612
rect 1590 588 1594 592
rect 1606 568 1610 572
rect 1566 548 1570 552
rect 1598 548 1602 552
rect 1414 538 1418 542
rect 1462 538 1466 542
rect 1470 538 1474 542
rect 1510 538 1514 542
rect 1542 538 1546 542
rect 1558 538 1562 542
rect 1438 528 1442 532
rect 1454 528 1458 532
rect 1478 528 1482 532
rect 1502 528 1506 532
rect 1550 528 1554 532
rect 1582 518 1586 522
rect 1446 508 1450 512
rect 1518 498 1522 502
rect 1462 488 1466 492
rect 1486 488 1490 492
rect 1422 468 1426 472
rect 1430 458 1434 462
rect 1438 458 1442 462
rect 1414 448 1418 452
rect 1446 428 1450 432
rect 1638 648 1642 652
rect 1662 648 1666 652
rect 1630 638 1634 642
rect 1622 598 1626 602
rect 1622 548 1626 552
rect 1654 598 1658 602
rect 1638 558 1642 562
rect 1638 538 1642 542
rect 1622 528 1626 532
rect 1646 528 1650 532
rect 1606 518 1610 522
rect 1606 488 1610 492
rect 1590 478 1594 482
rect 1510 448 1514 452
rect 1470 438 1474 442
rect 1478 418 1482 422
rect 1462 398 1466 402
rect 1446 378 1450 382
rect 1478 388 1482 392
rect 1462 358 1466 362
rect 1470 358 1474 362
rect 1398 338 1402 342
rect 1422 338 1426 342
rect 1302 328 1306 332
rect 1318 328 1322 332
rect 1382 328 1386 332
rect 1326 318 1330 322
rect 1238 308 1242 312
rect 1294 308 1298 312
rect 1302 308 1306 312
rect 1334 308 1338 312
rect 1358 308 1362 312
rect 1270 298 1274 302
rect 1254 288 1258 292
rect 1214 258 1218 262
rect 1182 248 1186 252
rect 1142 238 1146 242
rect 1174 238 1178 242
rect 1198 238 1202 242
rect 1134 198 1138 202
rect 1118 168 1122 172
rect 1134 158 1138 162
rect 814 128 818 132
rect 850 103 854 107
rect 857 103 861 107
rect 886 98 890 102
rect 918 98 922 102
rect 902 78 906 82
rect 966 138 970 142
rect 1110 148 1114 152
rect 1214 218 1218 222
rect 1158 188 1162 192
rect 1142 138 1146 142
rect 1198 158 1202 162
rect 1214 158 1218 162
rect 1318 288 1322 292
rect 1398 248 1402 252
rect 1362 203 1366 207
rect 1369 203 1373 207
rect 1278 178 1282 182
rect 1262 168 1266 172
rect 1270 168 1274 172
rect 1182 148 1186 152
rect 1230 148 1234 152
rect 1238 148 1242 152
rect 1174 138 1178 142
rect 1206 138 1210 142
rect 1214 138 1218 142
rect 1014 128 1018 132
rect 1078 128 1082 132
rect 1214 128 1218 132
rect 1118 88 1122 92
rect 1102 78 1106 82
rect 958 58 962 62
rect 1046 58 1050 62
rect 1158 58 1162 62
rect 726 8 730 12
rect 766 8 770 12
rect 782 8 786 12
rect 1102 8 1106 12
rect 1214 8 1218 12
rect 1230 8 1234 12
rect 1262 138 1266 142
rect 1302 158 1306 162
rect 1278 118 1282 122
rect 1254 108 1258 112
rect 1366 148 1370 152
rect 1422 148 1426 152
rect 1382 118 1386 122
rect 1318 108 1322 112
rect 1318 88 1322 92
rect 1246 58 1250 62
rect 1254 8 1258 12
rect 1278 8 1282 12
rect 1362 3 1366 7
rect 1369 3 1373 7
rect 1446 318 1450 322
rect 1502 408 1506 412
rect 1590 458 1594 462
rect 1526 448 1530 452
rect 1534 438 1538 442
rect 1518 358 1522 362
rect 1510 348 1514 352
rect 1526 348 1530 352
rect 1558 448 1562 452
rect 1542 358 1546 362
rect 1478 318 1482 322
rect 1550 348 1554 352
rect 1598 418 1602 422
rect 1574 348 1578 352
rect 1606 408 1610 412
rect 1622 398 1626 402
rect 1734 908 1738 912
rect 1718 878 1722 882
rect 1710 868 1714 872
rect 1782 888 1786 892
rect 1742 878 1746 882
rect 1774 878 1778 882
rect 1798 878 1802 882
rect 1782 868 1786 872
rect 1774 858 1778 862
rect 1718 848 1722 852
rect 1726 848 1730 852
rect 1750 848 1754 852
rect 1790 848 1794 852
rect 1806 848 1810 852
rect 1710 798 1714 802
rect 1718 798 1722 802
rect 1830 908 1834 912
rect 1830 898 1834 902
rect 1838 888 1842 892
rect 1966 928 1970 932
rect 1918 908 1922 912
rect 1882 903 1886 907
rect 1889 903 1893 907
rect 1870 898 1874 902
rect 1870 888 1874 892
rect 1902 888 1906 892
rect 1926 888 1930 892
rect 2070 908 2074 912
rect 1966 898 1970 902
rect 1966 888 1970 892
rect 1870 868 1874 872
rect 1942 868 1946 872
rect 1814 838 1818 842
rect 1782 828 1786 832
rect 1750 808 1754 812
rect 1734 768 1738 772
rect 1814 808 1818 812
rect 1878 848 1882 852
rect 1918 858 1922 862
rect 1934 848 1938 852
rect 1902 838 1906 842
rect 1894 818 1898 822
rect 1846 798 1850 802
rect 1862 798 1866 802
rect 1862 778 1866 782
rect 1798 758 1802 762
rect 1830 758 1834 762
rect 1758 748 1762 752
rect 1806 738 1810 742
rect 1742 728 1746 732
rect 1750 728 1754 732
rect 1758 718 1762 722
rect 1774 718 1778 722
rect 1718 698 1722 702
rect 1742 688 1746 692
rect 1726 678 1730 682
rect 1694 638 1698 642
rect 1694 598 1698 602
rect 1830 618 1834 622
rect 1750 588 1754 592
rect 1782 588 1786 592
rect 2198 998 2202 1002
rect 2174 948 2178 952
rect 2198 978 2202 982
rect 2190 958 2194 962
rect 2206 948 2210 952
rect 2206 928 2210 932
rect 2182 918 2186 922
rect 2118 908 2122 912
rect 2174 908 2178 912
rect 2310 1218 2314 1222
rect 2294 1168 2298 1172
rect 2326 1168 2330 1172
rect 2294 1158 2298 1162
rect 2318 1158 2322 1162
rect 2386 1203 2390 1207
rect 2393 1203 2397 1207
rect 2358 1158 2362 1162
rect 2366 1158 2370 1162
rect 2310 1148 2314 1152
rect 2342 1148 2346 1152
rect 2358 1148 2362 1152
rect 2318 1138 2322 1142
rect 2374 1138 2378 1142
rect 2390 1138 2394 1142
rect 2326 1128 2330 1132
rect 2358 1128 2362 1132
rect 2374 1128 2378 1132
rect 2310 1118 2314 1122
rect 2342 1118 2346 1122
rect 2262 1108 2266 1112
rect 2230 1068 2234 1072
rect 2286 1098 2290 1102
rect 2326 1088 2330 1092
rect 2342 1088 2346 1092
rect 2302 1078 2306 1082
rect 2350 1078 2354 1082
rect 2270 1068 2274 1072
rect 2222 1058 2226 1062
rect 2230 1028 2234 1032
rect 2222 978 2226 982
rect 2230 968 2234 972
rect 2366 1068 2370 1072
rect 2358 1058 2362 1062
rect 2262 1048 2266 1052
rect 2310 1048 2314 1052
rect 2294 978 2298 982
rect 2342 978 2346 982
rect 2270 958 2274 962
rect 2286 958 2290 962
rect 2342 958 2346 962
rect 2350 948 2354 952
rect 2366 1038 2370 1042
rect 2398 1128 2402 1132
rect 2422 1358 2426 1362
rect 2446 1438 2450 1442
rect 2438 1348 2442 1352
rect 2526 1498 2530 1502
rect 2462 1478 2466 1482
rect 2582 1478 2586 1482
rect 2590 1478 2594 1482
rect 2606 1478 2610 1482
rect 2614 1478 2618 1482
rect 2470 1458 2474 1462
rect 2478 1448 2482 1452
rect 2462 1348 2466 1352
rect 2494 1468 2498 1472
rect 2510 1468 2514 1472
rect 2606 1468 2610 1472
rect 2494 1448 2498 1452
rect 2566 1458 2570 1462
rect 2534 1438 2538 1442
rect 2542 1438 2546 1442
rect 2486 1428 2490 1432
rect 2494 1358 2498 1362
rect 2558 1428 2562 1432
rect 2550 1408 2554 1412
rect 2558 1398 2562 1402
rect 2566 1368 2570 1372
rect 2526 1348 2530 1352
rect 2550 1348 2554 1352
rect 2558 1348 2562 1352
rect 2582 1348 2586 1352
rect 2510 1338 2514 1342
rect 2462 1318 2466 1322
rect 2478 1318 2482 1322
rect 2438 1298 2442 1302
rect 2454 1298 2458 1302
rect 2430 1268 2434 1272
rect 2574 1338 2578 1342
rect 2518 1328 2522 1332
rect 2542 1328 2546 1332
rect 2534 1318 2538 1322
rect 2478 1308 2482 1312
rect 2494 1308 2498 1312
rect 2574 1328 2578 1332
rect 2494 1278 2498 1282
rect 2542 1278 2546 1282
rect 2558 1278 2562 1282
rect 2486 1268 2490 1272
rect 2446 1258 2450 1262
rect 2422 1238 2426 1242
rect 2414 1208 2418 1212
rect 2454 1208 2458 1212
rect 2462 1168 2466 1172
rect 2470 1158 2474 1162
rect 2526 1258 2530 1262
rect 2494 1208 2498 1212
rect 2510 1208 2514 1212
rect 2518 1188 2522 1192
rect 2494 1168 2498 1172
rect 2510 1158 2514 1162
rect 2446 1148 2450 1152
rect 2462 1148 2466 1152
rect 2430 1128 2434 1132
rect 2478 1128 2482 1132
rect 2454 1118 2458 1122
rect 2478 1118 2482 1122
rect 2446 1088 2450 1092
rect 2454 1088 2458 1092
rect 2406 1078 2410 1082
rect 2414 1078 2418 1082
rect 2454 1068 2458 1072
rect 2550 1158 2554 1162
rect 2494 1128 2498 1132
rect 2510 1128 2514 1132
rect 2526 1118 2530 1122
rect 2494 1078 2498 1082
rect 2518 1078 2522 1082
rect 2422 1058 2426 1062
rect 2366 1008 2370 1012
rect 2262 938 2266 942
rect 2278 938 2282 942
rect 2302 938 2306 942
rect 2310 938 2314 942
rect 2334 938 2338 942
rect 2222 928 2226 932
rect 2238 918 2242 922
rect 2254 908 2258 912
rect 2230 898 2234 902
rect 2350 928 2354 932
rect 2358 928 2362 932
rect 2294 908 2298 912
rect 2318 908 2322 912
rect 2262 888 2266 892
rect 2230 878 2234 882
rect 2110 868 2114 872
rect 2174 868 2178 872
rect 2310 888 2314 892
rect 2054 858 2058 862
rect 2142 858 2146 862
rect 1998 848 2002 852
rect 2038 848 2042 852
rect 1942 838 1946 842
rect 1950 838 1954 842
rect 2126 838 2130 842
rect 2062 818 2066 822
rect 1934 808 1938 812
rect 1886 768 1890 772
rect 1910 768 1914 772
rect 1882 703 1886 707
rect 1889 703 1893 707
rect 1886 688 1890 692
rect 1862 668 1866 672
rect 1846 648 1850 652
rect 1886 648 1890 652
rect 1990 748 1994 752
rect 2054 748 2058 752
rect 1974 738 1978 742
rect 2078 768 2082 772
rect 2134 808 2138 812
rect 2206 808 2210 812
rect 2142 798 2146 802
rect 2094 748 2098 752
rect 2126 748 2130 752
rect 2174 778 2178 782
rect 2238 798 2242 802
rect 2214 778 2218 782
rect 2278 778 2282 782
rect 2294 768 2298 772
rect 2262 758 2266 762
rect 2230 748 2234 752
rect 2086 738 2090 742
rect 2118 738 2122 742
rect 2158 738 2162 742
rect 2174 738 2178 742
rect 2286 738 2290 742
rect 2078 728 2082 732
rect 2198 728 2202 732
rect 1966 688 1970 692
rect 2062 688 2066 692
rect 1942 678 1946 682
rect 1974 678 1978 682
rect 1982 678 1986 682
rect 2046 678 2050 682
rect 1926 668 1930 672
rect 2022 668 2026 672
rect 2054 668 2058 672
rect 1950 658 1954 662
rect 1966 658 1970 662
rect 1990 658 1994 662
rect 1934 648 1938 652
rect 1974 648 1978 652
rect 1990 648 1994 652
rect 1854 638 1858 642
rect 1910 638 1914 642
rect 1950 638 1954 642
rect 1886 628 1890 632
rect 1838 558 1842 562
rect 1694 548 1698 552
rect 1886 548 1890 552
rect 1686 538 1690 542
rect 1710 538 1714 542
rect 1686 508 1690 512
rect 1686 498 1690 502
rect 1918 538 1922 542
rect 1750 528 1754 532
rect 1806 528 1810 532
rect 1942 528 1946 532
rect 1790 518 1794 522
rect 1750 508 1754 512
rect 1882 503 1886 507
rect 1889 503 1893 507
rect 1782 498 1786 502
rect 1734 488 1738 492
rect 1758 488 1762 492
rect 1862 488 1866 492
rect 1918 488 1922 492
rect 2030 658 2034 662
rect 2094 658 2098 662
rect 2014 648 2018 652
rect 2054 638 2058 642
rect 2006 628 2010 632
rect 2086 608 2090 612
rect 2062 588 2066 592
rect 2086 588 2090 592
rect 1982 518 1986 522
rect 1974 488 1978 492
rect 1670 478 1674 482
rect 1782 478 1786 482
rect 1814 478 1818 482
rect 1718 448 1722 452
rect 1782 458 1786 462
rect 1734 428 1738 432
rect 1742 428 1746 432
rect 1670 418 1674 422
rect 1702 398 1706 402
rect 1638 378 1642 382
rect 1654 378 1658 382
rect 1822 468 1826 472
rect 1846 468 1850 472
rect 1814 458 1818 462
rect 1838 458 1842 462
rect 1854 458 1858 462
rect 1894 468 1898 472
rect 1934 468 1938 472
rect 1886 458 1890 462
rect 1886 438 1890 442
rect 1846 428 1850 432
rect 1790 398 1794 402
rect 1742 368 1746 372
rect 1686 358 1690 362
rect 1822 398 1826 402
rect 1830 358 1834 362
rect 1654 348 1658 352
rect 1726 348 1730 352
rect 1798 348 1802 352
rect 1662 338 1666 342
rect 1742 338 1746 342
rect 1830 338 1834 342
rect 1582 328 1586 332
rect 1694 328 1698 332
rect 1542 308 1546 312
rect 1550 308 1554 312
rect 1526 288 1530 292
rect 1566 288 1570 292
rect 1574 288 1578 292
rect 1630 288 1634 292
rect 1502 278 1506 282
rect 1518 278 1522 282
rect 1534 278 1538 282
rect 1510 268 1514 272
rect 1582 268 1586 272
rect 1598 268 1602 272
rect 1622 268 1626 272
rect 1654 278 1658 282
rect 1686 268 1690 272
rect 1462 248 1466 252
rect 1534 248 1538 252
rect 1542 248 1546 252
rect 1630 248 1634 252
rect 1638 248 1642 252
rect 1494 238 1498 242
rect 1566 238 1570 242
rect 1614 238 1618 242
rect 1438 218 1442 222
rect 1582 218 1586 222
rect 1638 218 1642 222
rect 1454 188 1458 192
rect 1478 178 1482 182
rect 1566 158 1570 162
rect 1518 148 1522 152
rect 1462 128 1466 132
rect 1518 98 1522 102
rect 1670 248 1674 252
rect 1766 308 1770 312
rect 1830 308 1834 312
rect 1726 278 1730 282
rect 1758 268 1762 272
rect 1702 248 1706 252
rect 1718 248 1722 252
rect 1662 188 1666 192
rect 1654 178 1658 182
rect 1566 98 1570 102
rect 1614 88 1618 92
rect 1526 78 1530 82
rect 1566 78 1570 82
rect 1486 68 1490 72
rect 1526 68 1530 72
rect 1630 68 1634 72
rect 1798 278 1802 282
rect 1814 268 1818 272
rect 1742 248 1746 252
rect 1758 248 1762 252
rect 1774 248 1778 252
rect 1790 248 1794 252
rect 1870 378 1874 382
rect 1854 368 1858 372
rect 1910 448 1914 452
rect 1894 428 1898 432
rect 1902 388 1906 392
rect 1894 368 1898 372
rect 1862 348 1866 352
rect 1862 328 1866 332
rect 1882 303 1886 307
rect 1889 303 1893 307
rect 1870 298 1874 302
rect 1950 478 1954 482
rect 1982 468 1986 472
rect 1942 458 1946 462
rect 1934 408 1938 412
rect 1950 398 1954 402
rect 1934 368 1938 372
rect 1910 328 1914 332
rect 1918 328 1922 332
rect 1990 398 1994 402
rect 2118 688 2122 692
rect 2158 698 2162 702
rect 2198 698 2202 702
rect 2174 688 2178 692
rect 2126 658 2130 662
rect 2142 658 2146 662
rect 2134 638 2138 642
rect 2014 558 2018 562
rect 2022 558 2026 562
rect 2182 658 2186 662
rect 2190 648 2194 652
rect 2166 618 2170 622
rect 2134 608 2138 612
rect 2110 558 2114 562
rect 2166 558 2170 562
rect 2046 548 2050 552
rect 2078 538 2082 542
rect 2134 538 2138 542
rect 2062 528 2066 532
rect 2078 528 2082 532
rect 2118 528 2122 532
rect 2166 528 2170 532
rect 2142 518 2146 522
rect 2054 508 2058 512
rect 2070 488 2074 492
rect 2086 478 2090 482
rect 2142 468 2146 472
rect 2126 458 2130 462
rect 2014 448 2018 452
rect 1998 388 2002 392
rect 2126 398 2130 402
rect 2030 378 2034 382
rect 2102 378 2106 382
rect 2094 368 2098 372
rect 1982 358 1986 362
rect 2006 358 2010 362
rect 2030 358 2034 362
rect 2030 348 2034 352
rect 2086 348 2090 352
rect 2126 348 2130 352
rect 1974 338 1978 342
rect 1926 288 1930 292
rect 1958 328 1962 332
rect 1990 328 1994 332
rect 1990 318 1994 322
rect 1958 308 1962 312
rect 1974 278 1978 282
rect 1998 288 2002 292
rect 2030 338 2034 342
rect 2062 338 2066 342
rect 2078 338 2082 342
rect 2110 338 2114 342
rect 2030 328 2034 332
rect 2038 328 2042 332
rect 2030 278 2034 282
rect 2054 328 2058 332
rect 2102 328 2106 332
rect 2134 328 2138 332
rect 2046 308 2050 312
rect 2070 288 2074 292
rect 2118 288 2122 292
rect 2158 478 2162 482
rect 2166 478 2170 482
rect 2222 708 2226 712
rect 2198 608 2202 612
rect 2214 608 2218 612
rect 2206 538 2210 542
rect 2302 698 2306 702
rect 2278 688 2282 692
rect 2294 678 2298 682
rect 2254 668 2258 672
rect 2286 668 2290 672
rect 2358 898 2362 902
rect 2446 1048 2450 1052
rect 2430 1008 2434 1012
rect 2462 1008 2466 1012
rect 2386 1003 2390 1007
rect 2393 1003 2397 1007
rect 2470 978 2474 982
rect 2390 968 2394 972
rect 2382 958 2386 962
rect 2526 1068 2530 1072
rect 2542 1128 2546 1132
rect 2574 1268 2578 1272
rect 2566 1248 2570 1252
rect 2590 1168 2594 1172
rect 2614 1458 2618 1462
rect 2606 1438 2610 1442
rect 2630 1548 2634 1552
rect 2654 1568 2658 1572
rect 2718 1658 2722 1662
rect 2742 1728 2746 1732
rect 2894 1928 2898 1932
rect 2886 1918 2890 1922
rect 2846 1898 2850 1902
rect 2862 1898 2866 1902
rect 2822 1878 2826 1882
rect 2854 1878 2858 1882
rect 2774 1858 2778 1862
rect 2798 1848 2802 1852
rect 2814 1848 2818 1852
rect 2830 1848 2834 1852
rect 2766 1818 2770 1822
rect 2846 1858 2850 1862
rect 2806 1798 2810 1802
rect 2822 1798 2826 1802
rect 2838 1798 2842 1802
rect 2774 1758 2778 1762
rect 2878 1868 2882 1872
rect 2902 1918 2906 1922
rect 2906 1903 2910 1907
rect 2913 1903 2917 1907
rect 2990 2068 2994 2072
rect 3054 2128 3058 2132
rect 3062 2128 3066 2132
rect 3086 2128 3090 2132
rect 3046 2118 3050 2122
rect 2974 2048 2978 2052
rect 3030 2048 3034 2052
rect 3054 2068 3058 2072
rect 3046 2058 3050 2062
rect 3094 2088 3098 2092
rect 3150 2148 3154 2152
rect 3126 2108 3130 2112
rect 3134 2098 3138 2102
rect 3126 2088 3130 2092
rect 3158 2128 3162 2132
rect 3166 2098 3170 2102
rect 3158 2078 3162 2082
rect 3230 2328 3234 2332
rect 3246 2328 3250 2332
rect 3222 2318 3226 2322
rect 3222 2298 3226 2302
rect 3230 2298 3234 2302
rect 3230 2288 3234 2292
rect 3198 2268 3202 2272
rect 3230 2268 3234 2272
rect 3206 2258 3210 2262
rect 3222 2228 3226 2232
rect 3222 2218 3226 2222
rect 3198 2178 3202 2182
rect 3190 2158 3194 2162
rect 3214 2158 3218 2162
rect 3190 2148 3194 2152
rect 3230 2148 3234 2152
rect 3206 2138 3210 2142
rect 3198 2098 3202 2102
rect 3190 2078 3194 2082
rect 3110 2058 3114 2062
rect 3134 2058 3138 2062
rect 3086 2048 3090 2052
rect 3118 2048 3122 2052
rect 3006 2038 3010 2042
rect 3014 2038 3018 2042
rect 3038 2038 3042 2042
rect 3062 2038 3066 2042
rect 3086 2038 3090 2042
rect 2982 2018 2986 2022
rect 2998 1998 3002 2002
rect 2982 1958 2986 1962
rect 2974 1948 2978 1952
rect 3038 1948 3042 1952
rect 3046 1948 3050 1952
rect 3070 1948 3074 1952
rect 2958 1918 2962 1922
rect 2966 1918 2970 1922
rect 2950 1908 2954 1912
rect 2926 1878 2930 1882
rect 2990 1938 2994 1942
rect 3062 1938 3066 1942
rect 3078 1938 3082 1942
rect 2998 1928 3002 1932
rect 2958 1878 2962 1882
rect 2942 1868 2946 1872
rect 2982 1868 2986 1872
rect 2998 1868 3002 1872
rect 2878 1858 2882 1862
rect 2934 1848 2938 1852
rect 2942 1848 2946 1852
rect 2990 1848 2994 1852
rect 2950 1838 2954 1842
rect 2942 1788 2946 1792
rect 2886 1768 2890 1772
rect 2894 1768 2898 1772
rect 2854 1758 2858 1762
rect 2862 1758 2866 1762
rect 2798 1748 2802 1752
rect 2886 1758 2890 1762
rect 2918 1758 2922 1762
rect 2782 1738 2786 1742
rect 2790 1738 2794 1742
rect 2822 1738 2826 1742
rect 2878 1738 2882 1742
rect 2758 1708 2762 1712
rect 2766 1698 2770 1702
rect 2798 1698 2802 1702
rect 2870 1698 2874 1702
rect 2790 1678 2794 1682
rect 2958 1828 2962 1832
rect 2942 1738 2946 1742
rect 2950 1708 2954 1712
rect 2906 1703 2910 1707
rect 2913 1703 2917 1707
rect 2854 1678 2858 1682
rect 2870 1678 2874 1682
rect 2918 1678 2922 1682
rect 2926 1678 2930 1682
rect 2814 1668 2818 1672
rect 2830 1668 2834 1672
rect 2862 1668 2866 1672
rect 2782 1658 2786 1662
rect 2734 1648 2738 1652
rect 2750 1648 2754 1652
rect 2814 1648 2818 1652
rect 2822 1648 2826 1652
rect 2838 1648 2842 1652
rect 2870 1648 2874 1652
rect 2710 1618 2714 1622
rect 2734 1618 2738 1622
rect 2750 1598 2754 1602
rect 2766 1578 2770 1582
rect 2702 1568 2706 1572
rect 2646 1518 2650 1522
rect 2630 1466 2634 1470
rect 2622 1278 2626 1282
rect 2622 1258 2626 1262
rect 2614 1238 2618 1242
rect 2622 1218 2626 1222
rect 2614 1168 2618 1172
rect 2598 1158 2602 1162
rect 2710 1488 2714 1492
rect 2678 1478 2682 1482
rect 2670 1448 2674 1452
rect 2678 1448 2682 1452
rect 2878 1608 2882 1612
rect 2854 1568 2858 1572
rect 2870 1568 2874 1572
rect 2814 1558 2818 1562
rect 2846 1558 2850 1562
rect 2782 1528 2786 1532
rect 2782 1518 2786 1522
rect 2734 1508 2738 1512
rect 2750 1508 2754 1512
rect 2742 1498 2746 1502
rect 2750 1478 2754 1482
rect 2806 1508 2810 1512
rect 2910 1668 2914 1672
rect 2886 1598 2890 1602
rect 2894 1578 2898 1582
rect 2990 1838 2994 1842
rect 2982 1808 2986 1812
rect 2966 1748 2970 1752
rect 2974 1738 2978 1742
rect 2974 1718 2978 1722
rect 2974 1708 2978 1712
rect 2982 1688 2986 1692
rect 2974 1668 2978 1672
rect 2982 1668 2986 1672
rect 3038 1908 3042 1912
rect 3014 1898 3018 1902
rect 3046 1898 3050 1902
rect 3062 1898 3066 1902
rect 3102 2028 3106 2032
rect 3110 1938 3114 1942
rect 3102 1918 3106 1922
rect 3038 1878 3042 1882
rect 3046 1878 3050 1882
rect 3022 1858 3026 1862
rect 3006 1808 3010 1812
rect 3022 1798 3026 1802
rect 2998 1738 3002 1742
rect 3006 1738 3010 1742
rect 3070 1848 3074 1852
rect 3054 1808 3058 1812
rect 3110 1908 3114 1912
rect 3110 1878 3114 1882
rect 3094 1868 3098 1872
rect 3086 1838 3090 1842
rect 3078 1808 3082 1812
rect 3030 1758 3034 1762
rect 3078 1748 3082 1752
rect 3094 1748 3098 1752
rect 3158 1978 3162 1982
rect 3214 2128 3218 2132
rect 3230 2108 3234 2112
rect 3278 2438 3282 2442
rect 3294 2468 3298 2472
rect 3310 2408 3314 2412
rect 3294 2398 3298 2402
rect 3286 2388 3290 2392
rect 3302 2358 3306 2362
rect 3278 2338 3282 2342
rect 3294 2338 3298 2342
rect 3270 2328 3274 2332
rect 3270 2278 3274 2282
rect 3286 2278 3290 2282
rect 3262 2268 3266 2272
rect 3294 2258 3298 2262
rect 3246 2228 3250 2232
rect 3246 2168 3250 2172
rect 3270 2168 3274 2172
rect 3254 2158 3258 2162
rect 3262 2148 3266 2152
rect 3302 2158 3306 2162
rect 3294 2148 3298 2152
rect 3254 2138 3258 2142
rect 3246 2108 3250 2112
rect 3270 2098 3274 2102
rect 3238 2078 3242 2082
rect 3246 2068 3250 2072
rect 3230 2058 3234 2062
rect 3326 2488 3330 2492
rect 3422 2648 3426 2652
rect 3406 2628 3410 2632
rect 3410 2603 3414 2607
rect 3417 2603 3421 2607
rect 3438 2568 3442 2572
rect 3470 2648 3474 2652
rect 3494 2648 3498 2652
rect 3454 2618 3458 2622
rect 3478 2568 3482 2572
rect 3470 2558 3474 2562
rect 3622 2738 3626 2742
rect 3526 2728 3530 2732
rect 3614 2718 3618 2722
rect 3542 2708 3546 2712
rect 3542 2698 3546 2702
rect 3582 2698 3586 2702
rect 3526 2668 3530 2672
rect 3566 2688 3570 2692
rect 3590 2688 3594 2692
rect 3510 2648 3514 2652
rect 3534 2648 3538 2652
rect 3566 2648 3570 2652
rect 3566 2638 3570 2642
rect 3574 2638 3578 2642
rect 3590 2638 3594 2642
rect 3502 2628 3506 2632
rect 3502 2608 3506 2612
rect 3526 2588 3530 2592
rect 3526 2578 3530 2582
rect 3398 2548 3402 2552
rect 3494 2548 3498 2552
rect 3502 2548 3506 2552
rect 3518 2548 3522 2552
rect 3446 2538 3450 2542
rect 3646 2738 3650 2742
rect 3638 2718 3642 2722
rect 3630 2688 3634 2692
rect 3606 2668 3610 2672
rect 3630 2668 3634 2672
rect 3622 2648 3626 2652
rect 3710 2748 3714 2752
rect 3670 2738 3674 2742
rect 3758 2748 3762 2752
rect 3742 2728 3746 2732
rect 3774 2728 3778 2732
rect 3678 2718 3682 2722
rect 3750 2718 3754 2722
rect 3710 2708 3714 2712
rect 3670 2698 3674 2702
rect 3654 2678 3658 2682
rect 3694 2678 3698 2682
rect 3654 2658 3658 2662
rect 3710 2658 3714 2662
rect 3726 2658 3730 2662
rect 3654 2648 3658 2652
rect 3710 2648 3714 2652
rect 3590 2568 3594 2572
rect 3598 2568 3602 2572
rect 3614 2568 3618 2572
rect 3550 2558 3554 2562
rect 3606 2558 3610 2562
rect 3542 2548 3546 2552
rect 3398 2528 3402 2532
rect 3454 2528 3458 2532
rect 3494 2528 3498 2532
rect 3574 2518 3578 2522
rect 3398 2508 3402 2512
rect 3366 2488 3370 2492
rect 3382 2488 3386 2492
rect 3366 2478 3370 2482
rect 3390 2478 3394 2482
rect 3478 2508 3482 2512
rect 3438 2488 3442 2492
rect 3334 2468 3338 2472
rect 3374 2468 3378 2472
rect 3382 2468 3386 2472
rect 3406 2468 3410 2472
rect 3414 2458 3418 2462
rect 3334 2448 3338 2452
rect 3342 2448 3346 2452
rect 3326 2438 3330 2442
rect 3366 2448 3370 2452
rect 3398 2448 3402 2452
rect 3358 2428 3362 2432
rect 3414 2428 3418 2432
rect 3350 2368 3354 2372
rect 3342 2358 3346 2362
rect 3366 2418 3370 2422
rect 3342 2318 3346 2322
rect 3334 2268 3338 2272
rect 3326 2238 3330 2242
rect 3326 2228 3330 2232
rect 3358 2338 3362 2342
rect 3410 2403 3414 2407
rect 3417 2403 3421 2407
rect 3446 2468 3450 2472
rect 3470 2448 3474 2452
rect 3518 2478 3522 2482
rect 3542 2478 3546 2482
rect 3486 2468 3490 2472
rect 3494 2468 3498 2472
rect 3518 2468 3522 2472
rect 3502 2448 3506 2452
rect 3534 2448 3538 2452
rect 3558 2478 3562 2482
rect 3582 2478 3586 2482
rect 3670 2598 3674 2602
rect 3646 2578 3650 2582
rect 3638 2548 3642 2552
rect 3662 2548 3666 2552
rect 3726 2628 3730 2632
rect 3702 2578 3706 2582
rect 3694 2568 3698 2572
rect 3686 2558 3690 2562
rect 3614 2538 3618 2542
rect 3646 2538 3650 2542
rect 3678 2538 3682 2542
rect 3614 2468 3618 2472
rect 3574 2458 3578 2462
rect 3446 2438 3450 2442
rect 3510 2428 3514 2432
rect 3630 2508 3634 2512
rect 3758 2568 3762 2572
rect 3766 2548 3770 2552
rect 3742 2538 3746 2542
rect 3670 2508 3674 2512
rect 3718 2508 3722 2512
rect 3638 2498 3642 2502
rect 3654 2498 3658 2502
rect 3630 2448 3634 2452
rect 3622 2428 3626 2432
rect 3446 2368 3450 2372
rect 3462 2368 3466 2372
rect 3382 2348 3386 2352
rect 3366 2268 3370 2272
rect 3510 2348 3514 2352
rect 3454 2338 3458 2342
rect 3406 2328 3410 2332
rect 3422 2318 3426 2322
rect 3430 2278 3434 2282
rect 3454 2278 3458 2282
rect 3486 2278 3490 2282
rect 3398 2268 3402 2272
rect 3462 2268 3466 2272
rect 3478 2268 3482 2272
rect 3382 2258 3386 2262
rect 3454 2258 3458 2262
rect 3358 2248 3362 2252
rect 3374 2238 3378 2242
rect 3430 2238 3434 2242
rect 3334 2188 3338 2192
rect 3410 2203 3414 2207
rect 3417 2203 3421 2207
rect 3406 2188 3410 2192
rect 3398 2178 3402 2182
rect 3390 2168 3394 2172
rect 3478 2248 3482 2252
rect 3526 2388 3530 2392
rect 3550 2388 3554 2392
rect 3550 2378 3554 2382
rect 3598 2368 3602 2372
rect 3558 2348 3562 2352
rect 3598 2348 3602 2352
rect 3590 2338 3594 2342
rect 3622 2398 3626 2402
rect 3614 2378 3618 2382
rect 3614 2338 3618 2342
rect 3630 2338 3634 2342
rect 3542 2328 3546 2332
rect 3606 2328 3610 2332
rect 3542 2308 3546 2312
rect 3582 2308 3586 2312
rect 3590 2308 3594 2312
rect 3518 2298 3522 2302
rect 3518 2288 3522 2292
rect 3574 2288 3578 2292
rect 3574 2278 3578 2282
rect 3526 2268 3530 2272
rect 3534 2268 3538 2272
rect 3510 2258 3514 2262
rect 3510 2238 3514 2242
rect 3534 2248 3538 2252
rect 3518 2228 3522 2232
rect 3494 2218 3498 2222
rect 3510 2218 3514 2222
rect 3582 2258 3586 2262
rect 3606 2258 3610 2262
rect 3774 2508 3778 2512
rect 3734 2488 3738 2492
rect 3694 2478 3698 2482
rect 3702 2478 3706 2482
rect 3750 2478 3754 2482
rect 3646 2458 3650 2462
rect 3702 2458 3706 2462
rect 3694 2438 3698 2442
rect 3678 2418 3682 2422
rect 3662 2388 3666 2392
rect 3670 2388 3674 2392
rect 3702 2378 3706 2382
rect 3742 2398 3746 2402
rect 3662 2368 3666 2372
rect 3710 2368 3714 2372
rect 3734 2368 3738 2372
rect 3742 2358 3746 2362
rect 3686 2348 3690 2352
rect 3702 2348 3706 2352
rect 3638 2318 3642 2322
rect 3550 2248 3554 2252
rect 3558 2248 3562 2252
rect 3574 2238 3578 2242
rect 3454 2188 3458 2192
rect 3494 2188 3498 2192
rect 3550 2188 3554 2192
rect 3414 2158 3418 2162
rect 3430 2158 3434 2162
rect 3318 2148 3322 2152
rect 3350 2148 3354 2152
rect 3310 2138 3314 2142
rect 3310 2128 3314 2132
rect 3342 2128 3346 2132
rect 3342 2108 3346 2112
rect 3334 2098 3338 2102
rect 3302 2078 3306 2082
rect 3334 2078 3338 2082
rect 3238 2048 3242 2052
rect 3262 2048 3266 2052
rect 3190 2018 3194 2022
rect 3214 2008 3218 2012
rect 3150 1958 3154 1962
rect 3174 1958 3178 1962
rect 3150 1948 3154 1952
rect 3158 1938 3162 1942
rect 3174 1938 3178 1942
rect 3142 1928 3146 1932
rect 3126 1908 3130 1912
rect 3134 1888 3138 1892
rect 3286 2008 3290 2012
rect 3222 1988 3226 1992
rect 3262 1988 3266 1992
rect 3190 1928 3194 1932
rect 3158 1898 3162 1902
rect 3142 1868 3146 1872
rect 3150 1868 3154 1872
rect 3166 1868 3170 1872
rect 3238 1958 3242 1962
rect 3262 1958 3266 1962
rect 3270 1948 3274 1952
rect 3278 1938 3282 1942
rect 3302 2058 3306 2062
rect 3318 2058 3322 2062
rect 3310 2048 3314 2052
rect 3310 2018 3314 2022
rect 3294 1968 3298 1972
rect 3310 1958 3314 1962
rect 3326 1948 3330 1952
rect 3334 1948 3338 1952
rect 3302 1938 3306 1942
rect 3206 1908 3210 1912
rect 3214 1898 3218 1902
rect 3238 1908 3242 1912
rect 3230 1898 3234 1902
rect 3214 1888 3218 1892
rect 3158 1848 3162 1852
rect 3174 1848 3178 1852
rect 3190 1848 3194 1852
rect 3254 1908 3258 1912
rect 3254 1898 3258 1902
rect 3286 1898 3290 1902
rect 3246 1888 3250 1892
rect 3318 1928 3322 1932
rect 3326 1928 3330 1932
rect 3334 1908 3338 1912
rect 3238 1878 3242 1882
rect 3302 1878 3306 1882
rect 3310 1878 3314 1882
rect 3334 1878 3338 1882
rect 3278 1868 3282 1872
rect 3238 1858 3242 1862
rect 3270 1858 3274 1862
rect 3302 1858 3306 1862
rect 3334 1858 3338 1862
rect 3198 1838 3202 1842
rect 3214 1838 3218 1842
rect 3118 1828 3122 1832
rect 3118 1768 3122 1772
rect 3262 1848 3266 1852
rect 3278 1838 3282 1842
rect 3286 1838 3290 1842
rect 3222 1828 3226 1832
rect 3270 1818 3274 1822
rect 3238 1798 3242 1802
rect 3166 1768 3170 1772
rect 3190 1768 3194 1772
rect 3134 1758 3138 1762
rect 3126 1748 3130 1752
rect 3014 1678 3018 1682
rect 2998 1668 3002 1672
rect 3046 1718 3050 1722
rect 3062 1718 3066 1722
rect 3078 1708 3082 1712
rect 3046 1678 3050 1682
rect 3006 1658 3010 1662
rect 3030 1658 3034 1662
rect 2990 1608 2994 1612
rect 2942 1578 2946 1582
rect 2998 1578 3002 1582
rect 2918 1568 2922 1572
rect 2982 1568 2986 1572
rect 2886 1558 2890 1562
rect 2942 1558 2946 1562
rect 2966 1558 2970 1562
rect 2894 1548 2898 1552
rect 2910 1548 2914 1552
rect 2870 1538 2874 1542
rect 2854 1518 2858 1522
rect 2886 1508 2890 1512
rect 2846 1498 2850 1502
rect 2854 1498 2858 1502
rect 2814 1488 2818 1492
rect 2838 1488 2842 1492
rect 2758 1448 2762 1452
rect 2798 1448 2802 1452
rect 2654 1438 2658 1442
rect 2686 1438 2690 1442
rect 2718 1428 2722 1432
rect 2934 1538 2938 1542
rect 2998 1548 3002 1552
rect 2982 1538 2986 1542
rect 2974 1528 2978 1532
rect 2906 1503 2910 1507
rect 2913 1503 2917 1507
rect 2942 1458 2946 1462
rect 2758 1358 2762 1362
rect 2766 1358 2770 1362
rect 2646 1318 2650 1322
rect 2686 1318 2690 1322
rect 2686 1308 2690 1312
rect 2646 1298 2650 1302
rect 2726 1288 2730 1292
rect 2742 1278 2746 1282
rect 2846 1418 2850 1422
rect 2870 1418 2874 1422
rect 2894 1418 2898 1422
rect 2846 1408 2850 1412
rect 2790 1368 2794 1372
rect 2798 1358 2802 1362
rect 2854 1378 2858 1382
rect 2894 1378 2898 1382
rect 2814 1348 2818 1352
rect 2838 1338 2842 1342
rect 2798 1308 2802 1312
rect 2782 1298 2786 1302
rect 2814 1298 2818 1302
rect 2838 1318 2842 1322
rect 2830 1288 2834 1292
rect 2838 1288 2842 1292
rect 2830 1278 2834 1282
rect 2774 1268 2778 1272
rect 2646 1248 2650 1252
rect 2646 1198 2650 1202
rect 2822 1168 2826 1172
rect 2742 1158 2746 1162
rect 2630 1148 2634 1152
rect 2782 1148 2786 1152
rect 2566 1128 2570 1132
rect 2574 1128 2578 1132
rect 2606 1128 2610 1132
rect 2662 1128 2666 1132
rect 2590 1118 2594 1122
rect 2582 1108 2586 1112
rect 2558 1088 2562 1092
rect 2630 1118 2634 1122
rect 2638 1118 2642 1122
rect 2598 1108 2602 1112
rect 2606 1108 2610 1112
rect 2598 1088 2602 1092
rect 2542 1068 2546 1072
rect 2598 1068 2602 1072
rect 2606 1068 2610 1072
rect 2494 1058 2498 1062
rect 2534 1058 2538 1062
rect 2502 1048 2506 1052
rect 2494 968 2498 972
rect 2478 958 2482 962
rect 2422 948 2426 952
rect 2478 948 2482 952
rect 2502 948 2506 952
rect 2526 958 2530 962
rect 2534 948 2538 952
rect 2438 938 2442 942
rect 2478 938 2482 942
rect 2486 938 2490 942
rect 2510 938 2514 942
rect 2390 928 2394 932
rect 2454 928 2458 932
rect 2374 908 2378 912
rect 2342 878 2346 882
rect 2366 878 2370 882
rect 2326 818 2330 822
rect 2326 798 2330 802
rect 2406 888 2410 892
rect 2446 898 2450 902
rect 2438 888 2442 892
rect 2430 878 2434 882
rect 2534 928 2538 932
rect 2462 898 2466 902
rect 2486 898 2490 902
rect 2414 858 2418 862
rect 2382 838 2386 842
rect 2366 828 2370 832
rect 2386 803 2390 807
rect 2393 803 2397 807
rect 2374 798 2378 802
rect 2358 778 2362 782
rect 2334 768 2338 772
rect 2326 748 2330 752
rect 2318 688 2322 692
rect 2350 678 2354 682
rect 2518 908 2522 912
rect 2534 898 2538 902
rect 2478 878 2482 882
rect 2526 878 2530 882
rect 2486 868 2490 872
rect 2494 868 2498 872
rect 2454 858 2458 862
rect 2430 848 2434 852
rect 2462 848 2466 852
rect 2566 1058 2570 1062
rect 2582 1058 2586 1062
rect 2590 1038 2594 1042
rect 2558 968 2562 972
rect 2566 968 2570 972
rect 2582 958 2586 962
rect 2654 1088 2658 1092
rect 2638 1078 2642 1082
rect 2726 1118 2730 1122
rect 2774 1118 2778 1122
rect 2742 1098 2746 1102
rect 2678 1088 2682 1092
rect 2710 1078 2714 1082
rect 2758 1088 2762 1092
rect 2686 1068 2690 1072
rect 2718 1068 2722 1072
rect 2622 1058 2626 1062
rect 2646 1058 2650 1062
rect 2598 968 2602 972
rect 2694 1048 2698 1052
rect 2726 1048 2730 1052
rect 2734 1048 2738 1052
rect 2670 978 2674 982
rect 2646 958 2650 962
rect 2622 948 2626 952
rect 2654 948 2658 952
rect 2686 948 2690 952
rect 2582 938 2586 942
rect 2598 938 2602 942
rect 2646 938 2650 942
rect 2662 938 2666 942
rect 2614 928 2618 932
rect 2686 928 2690 932
rect 2558 908 2562 912
rect 2590 908 2594 912
rect 2558 898 2562 902
rect 2606 878 2610 882
rect 2510 838 2514 842
rect 2542 838 2546 842
rect 2422 828 2426 832
rect 2494 828 2498 832
rect 2462 808 2466 812
rect 2430 768 2434 772
rect 2454 768 2458 772
rect 2406 738 2410 742
rect 2422 738 2426 742
rect 2374 728 2378 732
rect 2406 728 2410 732
rect 2366 678 2370 682
rect 2438 728 2442 732
rect 2454 728 2458 732
rect 2446 698 2450 702
rect 2438 688 2442 692
rect 2446 688 2450 692
rect 2638 878 2642 882
rect 2686 878 2690 882
rect 2702 878 2706 882
rect 2582 868 2586 872
rect 2614 868 2618 872
rect 2630 868 2634 872
rect 2662 868 2666 872
rect 2670 868 2674 872
rect 2694 868 2698 872
rect 2622 858 2626 862
rect 2646 858 2650 862
rect 2678 858 2682 862
rect 2566 808 2570 812
rect 2550 798 2554 802
rect 2526 778 2530 782
rect 2614 808 2618 812
rect 2526 768 2530 772
rect 2582 768 2586 772
rect 2494 748 2498 752
rect 2510 748 2514 752
rect 2478 738 2482 742
rect 2494 738 2498 742
rect 2470 728 2474 732
rect 2486 728 2490 732
rect 2510 698 2514 702
rect 2470 678 2474 682
rect 2230 658 2234 662
rect 2246 658 2250 662
rect 2262 658 2266 662
rect 2334 658 2338 662
rect 2358 658 2362 662
rect 2406 658 2410 662
rect 2238 598 2242 602
rect 2238 558 2242 562
rect 2302 648 2306 652
rect 2310 648 2314 652
rect 2350 648 2354 652
rect 2254 618 2258 622
rect 2286 618 2290 622
rect 2270 608 2274 612
rect 2318 608 2322 612
rect 2326 598 2330 602
rect 2262 568 2266 572
rect 2254 558 2258 562
rect 2302 558 2306 562
rect 2246 548 2250 552
rect 2214 528 2218 532
rect 2214 508 2218 512
rect 2206 478 2210 482
rect 2182 458 2186 462
rect 2278 538 2282 542
rect 2294 518 2298 522
rect 2278 498 2282 502
rect 2222 458 2226 462
rect 2254 458 2258 462
rect 2262 458 2266 462
rect 2278 458 2282 462
rect 2214 428 2218 432
rect 2198 368 2202 372
rect 2158 288 2162 292
rect 2046 278 2050 282
rect 2062 278 2066 282
rect 2014 268 2018 272
rect 1878 258 1882 262
rect 1974 258 1978 262
rect 1814 248 1818 252
rect 1926 248 1930 252
rect 1934 248 1938 252
rect 1878 238 1882 242
rect 1982 238 1986 242
rect 1998 238 2002 242
rect 1806 228 1810 232
rect 1782 218 1786 222
rect 1734 198 1738 202
rect 1702 178 1706 182
rect 1702 158 1706 162
rect 1846 168 1850 172
rect 1814 148 1818 152
rect 1742 138 1746 142
rect 1758 118 1762 122
rect 1814 98 1818 102
rect 1830 98 1834 102
rect 1750 78 1754 82
rect 1694 48 1698 52
rect 1982 218 1986 222
rect 2038 228 2042 232
rect 2078 228 2082 232
rect 2006 208 2010 212
rect 2014 208 2018 212
rect 1902 188 1906 192
rect 1894 128 1898 132
rect 1882 103 1886 107
rect 1889 103 1893 107
rect 1918 178 1922 182
rect 2102 278 2106 282
rect 2110 278 2114 282
rect 2094 248 2098 252
rect 2086 158 2090 162
rect 1926 148 1930 152
rect 1982 148 1986 152
rect 2118 168 2122 172
rect 2102 158 2106 162
rect 2214 318 2218 322
rect 2214 288 2218 292
rect 2198 278 2202 282
rect 2206 278 2210 282
rect 2150 248 2154 252
rect 2158 248 2162 252
rect 2166 248 2170 252
rect 2182 238 2186 242
rect 2198 248 2202 252
rect 2206 248 2210 252
rect 2166 208 2170 212
rect 2190 208 2194 212
rect 2270 438 2274 442
rect 2230 428 2234 432
rect 2238 378 2242 382
rect 2246 368 2250 372
rect 2230 358 2234 362
rect 2238 348 2242 352
rect 2270 348 2274 352
rect 2286 348 2290 352
rect 2238 278 2242 282
rect 2246 278 2250 282
rect 2386 603 2390 607
rect 2393 603 2397 607
rect 2438 598 2442 602
rect 2486 668 2490 672
rect 2470 648 2474 652
rect 2502 648 2506 652
rect 2566 748 2570 752
rect 2814 1128 2818 1132
rect 2814 1108 2818 1112
rect 2782 1088 2786 1092
rect 2854 1358 2858 1362
rect 2870 1358 2874 1362
rect 2886 1358 2890 1362
rect 2862 1348 2866 1352
rect 2870 1338 2874 1342
rect 2846 1268 2850 1272
rect 2846 1258 2850 1262
rect 2854 1238 2858 1242
rect 2838 1228 2842 1232
rect 2838 1198 2842 1202
rect 2886 1308 2890 1312
rect 2878 1248 2882 1252
rect 2862 1188 2866 1192
rect 2854 1178 2858 1182
rect 2846 1158 2850 1162
rect 2830 1078 2834 1082
rect 2838 1078 2842 1082
rect 2862 1158 2866 1162
rect 2870 1148 2874 1152
rect 2902 1348 2906 1352
rect 2906 1303 2910 1307
rect 2913 1303 2917 1307
rect 2902 1268 2906 1272
rect 2910 1258 2914 1262
rect 2902 1158 2906 1162
rect 2894 1138 2898 1142
rect 2862 1128 2866 1132
rect 2870 1128 2874 1132
rect 2862 1078 2866 1082
rect 2798 1058 2802 1062
rect 2814 1058 2818 1062
rect 2838 1058 2842 1062
rect 2766 1048 2770 1052
rect 2790 1048 2794 1052
rect 2806 1048 2810 1052
rect 2758 1038 2762 1042
rect 2750 1008 2754 1012
rect 2726 998 2730 1002
rect 2742 998 2746 1002
rect 2774 998 2778 1002
rect 2718 958 2722 962
rect 2790 988 2794 992
rect 2782 968 2786 972
rect 2734 948 2738 952
rect 2750 878 2754 882
rect 2734 868 2738 872
rect 2702 838 2706 842
rect 2654 828 2658 832
rect 2662 818 2666 822
rect 2694 808 2698 812
rect 2766 908 2770 912
rect 2766 878 2770 882
rect 2838 958 2842 962
rect 2814 948 2818 952
rect 2806 938 2810 942
rect 2798 928 2802 932
rect 2846 948 2850 952
rect 2838 938 2842 942
rect 2862 1038 2866 1042
rect 2906 1103 2910 1107
rect 2913 1103 2917 1107
rect 2918 1058 2922 1062
rect 3094 1718 3098 1722
rect 3094 1678 3098 1682
rect 3102 1678 3106 1682
rect 3038 1638 3042 1642
rect 3022 1618 3026 1622
rect 3014 1568 3018 1572
rect 3086 1658 3090 1662
rect 3054 1608 3058 1612
rect 3070 1608 3074 1612
rect 3030 1568 3034 1572
rect 3070 1598 3074 1602
rect 3054 1558 3058 1562
rect 3038 1548 3042 1552
rect 3094 1588 3098 1592
rect 3086 1548 3090 1552
rect 3078 1538 3082 1542
rect 3126 1728 3130 1732
rect 3142 1728 3146 1732
rect 3134 1688 3138 1692
rect 3158 1748 3162 1752
rect 3174 1748 3178 1752
rect 3222 1748 3226 1752
rect 3206 1718 3210 1722
rect 3206 1698 3210 1702
rect 3318 1798 3322 1802
rect 3294 1778 3298 1782
rect 3366 2118 3370 2122
rect 3358 2068 3362 2072
rect 3358 2048 3362 2052
rect 3382 2068 3386 2072
rect 3390 2058 3394 2062
rect 3526 2168 3530 2172
rect 3478 2148 3482 2152
rect 3502 2148 3506 2152
rect 3422 2128 3426 2132
rect 3438 2098 3442 2102
rect 3438 2078 3442 2082
rect 3470 2138 3474 2142
rect 3454 2078 3458 2082
rect 3446 2068 3450 2072
rect 3438 2058 3442 2062
rect 3382 2048 3386 2052
rect 3398 2048 3402 2052
rect 3470 2048 3474 2052
rect 3502 2098 3506 2102
rect 3478 2038 3482 2042
rect 3374 2028 3378 2032
rect 3414 2028 3418 2032
rect 3462 2028 3466 2032
rect 3566 2178 3570 2182
rect 3670 2328 3674 2332
rect 3654 2308 3658 2312
rect 3678 2298 3682 2302
rect 3646 2288 3650 2292
rect 3686 2278 3690 2282
rect 3710 2268 3714 2272
rect 3686 2258 3690 2262
rect 3694 2248 3698 2252
rect 3654 2238 3658 2242
rect 3606 2218 3610 2222
rect 3654 2218 3658 2222
rect 3670 2218 3674 2222
rect 3590 2188 3594 2192
rect 3582 2178 3586 2182
rect 3598 2178 3602 2182
rect 3662 2178 3666 2182
rect 3558 2158 3562 2162
rect 3574 2158 3578 2162
rect 3606 2158 3610 2162
rect 3526 2128 3530 2132
rect 3542 2048 3546 2052
rect 3510 2038 3514 2042
rect 3486 2018 3490 2022
rect 3398 2008 3402 2012
rect 3486 2008 3490 2012
rect 3410 2003 3414 2007
rect 3417 2003 3421 2007
rect 3526 2038 3530 2042
rect 3550 2038 3554 2042
rect 3566 2148 3570 2152
rect 3606 2088 3610 2092
rect 3574 2078 3578 2082
rect 3590 2068 3594 2072
rect 3566 2058 3570 2062
rect 3582 2058 3586 2062
rect 3734 2348 3738 2352
rect 3742 2338 3746 2342
rect 3734 2278 3738 2282
rect 3766 2258 3770 2262
rect 3734 2248 3738 2252
rect 3750 2248 3754 2252
rect 3718 2238 3722 2242
rect 3758 2238 3762 2242
rect 3726 2228 3730 2232
rect 3678 2158 3682 2162
rect 3638 2148 3642 2152
rect 3710 2168 3714 2172
rect 3718 2168 3722 2172
rect 3726 2158 3730 2162
rect 3654 2128 3658 2132
rect 3686 2128 3690 2132
rect 3678 2118 3682 2122
rect 3694 2118 3698 2122
rect 3678 2108 3682 2112
rect 3638 2088 3642 2092
rect 3630 2068 3634 2072
rect 3574 2018 3578 2022
rect 3526 2008 3530 2012
rect 3398 1958 3402 1962
rect 3446 1958 3450 1962
rect 3478 1958 3482 1962
rect 3510 1958 3514 1962
rect 3518 1958 3522 1962
rect 3374 1938 3378 1942
rect 3542 1998 3546 2002
rect 3638 2038 3642 2042
rect 3638 2028 3642 2032
rect 3622 1998 3626 2002
rect 3614 1988 3618 1992
rect 3534 1968 3538 1972
rect 3590 1968 3594 1972
rect 3606 1968 3610 1972
rect 3470 1948 3474 1952
rect 3406 1938 3410 1942
rect 3462 1938 3466 1942
rect 3486 1938 3490 1942
rect 3422 1918 3426 1922
rect 3382 1908 3386 1912
rect 3366 1898 3370 1902
rect 3390 1898 3394 1902
rect 3374 1848 3378 1852
rect 3382 1838 3386 1842
rect 3310 1768 3314 1772
rect 3350 1768 3354 1772
rect 3302 1758 3306 1762
rect 3286 1748 3290 1752
rect 3246 1738 3250 1742
rect 3222 1708 3226 1712
rect 3294 1738 3298 1742
rect 3254 1708 3258 1712
rect 3262 1698 3266 1702
rect 3158 1688 3162 1692
rect 3246 1688 3250 1692
rect 3142 1678 3146 1682
rect 3222 1678 3226 1682
rect 3166 1668 3170 1672
rect 3118 1648 3122 1652
rect 3110 1578 3114 1582
rect 3166 1648 3170 1652
rect 3182 1648 3186 1652
rect 3198 1608 3202 1612
rect 3174 1598 3178 1602
rect 3166 1588 3170 1592
rect 3214 1588 3218 1592
rect 3134 1578 3138 1582
rect 3110 1568 3114 1572
rect 3118 1568 3122 1572
rect 3190 1568 3194 1572
rect 3118 1558 3122 1562
rect 3038 1528 3042 1532
rect 3102 1528 3106 1532
rect 3030 1488 3034 1492
rect 2958 1468 2962 1472
rect 2998 1468 3002 1472
rect 3046 1518 3050 1522
rect 3094 1498 3098 1502
rect 2966 1458 2970 1462
rect 3006 1458 3010 1462
rect 2982 1448 2986 1452
rect 2950 1408 2954 1412
rect 3038 1408 3042 1412
rect 3046 1388 3050 1392
rect 3022 1378 3026 1382
rect 2974 1368 2978 1372
rect 3014 1368 3018 1372
rect 2966 1358 2970 1362
rect 2998 1358 3002 1362
rect 3022 1358 3026 1362
rect 2942 1328 2946 1332
rect 2958 1328 2962 1332
rect 3006 1348 3010 1352
rect 3030 1348 3034 1352
rect 3022 1338 3026 1342
rect 3014 1328 3018 1332
rect 2990 1318 2994 1322
rect 2934 1308 2938 1312
rect 2966 1308 2970 1312
rect 2998 1308 3002 1312
rect 2974 1298 2978 1302
rect 2974 1288 2978 1292
rect 2950 1278 2954 1282
rect 2934 1248 2938 1252
rect 2982 1278 2986 1282
rect 2950 1258 2954 1262
rect 2974 1248 2978 1252
rect 2958 1208 2962 1212
rect 2974 1208 2978 1212
rect 2942 1198 2946 1202
rect 2950 1198 2954 1202
rect 2942 1188 2946 1192
rect 2950 1168 2954 1172
rect 2958 1158 2962 1162
rect 2958 1148 2962 1152
rect 2966 1128 2970 1132
rect 2934 1108 2938 1112
rect 2942 1088 2946 1092
rect 2982 1198 2986 1202
rect 2990 1158 2994 1162
rect 3006 1298 3010 1302
rect 3014 1278 3018 1282
rect 3030 1328 3034 1332
rect 3238 1668 3242 1672
rect 3358 1758 3362 1762
rect 3422 1878 3426 1882
rect 3574 1958 3578 1962
rect 3558 1948 3562 1952
rect 3606 1948 3610 1952
rect 3550 1938 3554 1942
rect 3566 1938 3570 1942
rect 3606 1938 3610 1942
rect 3638 1998 3642 2002
rect 3630 1968 3634 1972
rect 3670 2058 3674 2062
rect 3670 2038 3674 2042
rect 3686 2028 3690 2032
rect 3662 2008 3666 2012
rect 3646 1978 3650 1982
rect 3734 2138 3738 2142
rect 3726 2098 3730 2102
rect 3718 2088 3722 2092
rect 3718 2078 3722 2082
rect 3710 2058 3714 2062
rect 3742 2088 3746 2092
rect 3734 2078 3738 2082
rect 3742 2068 3746 2072
rect 3726 2038 3730 2042
rect 3742 2038 3746 2042
rect 3742 2018 3746 2022
rect 3774 2108 3778 2112
rect 3766 2088 3770 2092
rect 3758 1998 3762 2002
rect 3702 1968 3706 1972
rect 3734 1968 3738 1972
rect 3638 1948 3642 1952
rect 3662 1948 3666 1952
rect 3670 1948 3674 1952
rect 3654 1938 3658 1942
rect 3446 1928 3450 1932
rect 3502 1928 3506 1932
rect 3526 1928 3530 1932
rect 3558 1928 3562 1932
rect 3582 1928 3586 1932
rect 3630 1928 3634 1932
rect 3662 1928 3666 1932
rect 3454 1908 3458 1912
rect 3446 1898 3450 1902
rect 3534 1888 3538 1892
rect 3470 1878 3474 1882
rect 3502 1878 3506 1882
rect 3574 1878 3578 1882
rect 3438 1868 3442 1872
rect 3478 1868 3482 1872
rect 3486 1868 3490 1872
rect 3502 1868 3506 1872
rect 3398 1828 3402 1832
rect 3410 1803 3414 1807
rect 3417 1803 3421 1807
rect 3470 1858 3474 1862
rect 3590 1888 3594 1892
rect 3662 1898 3666 1902
rect 3598 1878 3602 1882
rect 3622 1878 3626 1882
rect 3638 1878 3642 1882
rect 3606 1868 3610 1872
rect 3542 1858 3546 1862
rect 3582 1858 3586 1862
rect 3446 1838 3450 1842
rect 3494 1848 3498 1852
rect 3510 1848 3514 1852
rect 3534 1848 3538 1852
rect 3558 1838 3562 1842
rect 3582 1838 3586 1842
rect 3638 1868 3642 1872
rect 3654 1868 3658 1872
rect 3630 1848 3634 1852
rect 3694 1888 3698 1892
rect 3686 1878 3690 1882
rect 3694 1868 3698 1872
rect 3726 1878 3730 1882
rect 3726 1868 3730 1872
rect 3742 1938 3746 1942
rect 3670 1838 3674 1842
rect 3710 1838 3714 1842
rect 3486 1828 3490 1832
rect 3542 1828 3546 1832
rect 3614 1828 3618 1832
rect 3670 1828 3674 1832
rect 3702 1828 3706 1832
rect 3470 1808 3474 1812
rect 3470 1768 3474 1772
rect 3718 1818 3722 1822
rect 3502 1808 3506 1812
rect 3566 1798 3570 1802
rect 3510 1788 3514 1792
rect 3550 1788 3554 1792
rect 3518 1768 3522 1772
rect 3526 1768 3530 1772
rect 3606 1768 3610 1772
rect 3638 1768 3642 1772
rect 3542 1758 3546 1762
rect 3558 1758 3562 1762
rect 3590 1758 3594 1762
rect 3606 1758 3610 1762
rect 3406 1748 3410 1752
rect 3446 1748 3450 1752
rect 3486 1748 3490 1752
rect 3318 1738 3322 1742
rect 3342 1738 3346 1742
rect 3326 1698 3330 1702
rect 3374 1718 3378 1722
rect 3334 1678 3338 1682
rect 3478 1728 3482 1732
rect 3390 1678 3394 1682
rect 3286 1668 3290 1672
rect 3310 1668 3314 1672
rect 3326 1668 3330 1672
rect 3366 1668 3370 1672
rect 3390 1668 3394 1672
rect 3414 1668 3418 1672
rect 3254 1648 3258 1652
rect 3262 1648 3266 1652
rect 3230 1638 3234 1642
rect 3254 1558 3258 1562
rect 3134 1548 3138 1552
rect 3150 1548 3154 1552
rect 3222 1548 3226 1552
rect 3134 1528 3138 1532
rect 3118 1478 3122 1482
rect 3062 1468 3066 1472
rect 3214 1538 3218 1542
rect 3238 1538 3242 1542
rect 3166 1528 3170 1532
rect 3390 1648 3394 1652
rect 3462 1708 3466 1712
rect 3486 1678 3490 1682
rect 3430 1658 3434 1662
rect 3462 1658 3466 1662
rect 3334 1638 3338 1642
rect 3358 1638 3362 1642
rect 3422 1638 3426 1642
rect 3462 1638 3466 1642
rect 3486 1638 3490 1642
rect 3294 1588 3298 1592
rect 3278 1558 3282 1562
rect 3286 1558 3290 1562
rect 3238 1528 3242 1532
rect 3270 1528 3274 1532
rect 3222 1518 3226 1522
rect 3230 1508 3234 1512
rect 3150 1498 3154 1502
rect 3182 1498 3186 1502
rect 3190 1498 3194 1502
rect 3174 1488 3178 1492
rect 3166 1478 3170 1482
rect 3214 1478 3218 1482
rect 3158 1468 3162 1472
rect 3126 1458 3130 1462
rect 3078 1448 3082 1452
rect 3086 1418 3090 1422
rect 3054 1358 3058 1362
rect 3054 1348 3058 1352
rect 3062 1338 3066 1342
rect 3046 1268 3050 1272
rect 2982 1148 2986 1152
rect 3118 1388 3122 1392
rect 3126 1378 3130 1382
rect 3110 1348 3114 1352
rect 3150 1398 3154 1402
rect 3142 1368 3146 1372
rect 3166 1378 3170 1382
rect 3086 1318 3090 1322
rect 3142 1338 3146 1342
rect 3102 1328 3106 1332
rect 3070 1288 3074 1292
rect 3094 1288 3098 1292
rect 3062 1258 3066 1262
rect 3022 1208 3026 1212
rect 3062 1188 3066 1192
rect 3062 1168 3066 1172
rect 3142 1318 3146 1322
rect 3182 1338 3186 1342
rect 3214 1468 3218 1472
rect 3254 1518 3258 1522
rect 3246 1478 3250 1482
rect 3238 1458 3242 1462
rect 3254 1458 3258 1462
rect 3262 1458 3266 1462
rect 3222 1448 3226 1452
rect 3198 1418 3202 1422
rect 3214 1358 3218 1362
rect 3198 1348 3202 1352
rect 3174 1308 3178 1312
rect 3134 1298 3138 1302
rect 3166 1298 3170 1302
rect 3110 1278 3114 1282
rect 3102 1248 3106 1252
rect 3094 1238 3098 1242
rect 3102 1218 3106 1222
rect 3078 1208 3082 1212
rect 3070 1158 3074 1162
rect 3142 1278 3146 1282
rect 3134 1268 3138 1272
rect 3238 1408 3242 1412
rect 3230 1348 3234 1352
rect 3254 1368 3258 1372
rect 3254 1348 3258 1352
rect 3230 1318 3234 1322
rect 3222 1308 3226 1312
rect 3190 1298 3194 1302
rect 3230 1298 3234 1302
rect 3214 1288 3218 1292
rect 3238 1278 3242 1282
rect 3410 1603 3414 1607
rect 3417 1603 3421 1607
rect 3454 1588 3458 1592
rect 3366 1578 3370 1582
rect 3398 1578 3402 1582
rect 3310 1568 3314 1572
rect 3318 1558 3322 1562
rect 3358 1558 3362 1562
rect 3286 1538 3290 1542
rect 3390 1568 3394 1572
rect 3422 1568 3426 1572
rect 3374 1548 3378 1552
rect 3350 1538 3354 1542
rect 3398 1538 3402 1542
rect 3414 1538 3418 1542
rect 3310 1528 3314 1532
rect 3318 1528 3322 1532
rect 3302 1518 3306 1522
rect 3286 1508 3290 1512
rect 3294 1508 3298 1512
rect 3318 1508 3322 1512
rect 3294 1468 3298 1472
rect 3294 1418 3298 1422
rect 3294 1358 3298 1362
rect 3278 1328 3282 1332
rect 3302 1328 3306 1332
rect 3286 1288 3290 1292
rect 3342 1518 3346 1522
rect 3342 1508 3346 1512
rect 3326 1498 3330 1502
rect 3366 1468 3370 1472
rect 3358 1448 3362 1452
rect 3326 1438 3330 1442
rect 3334 1428 3338 1432
rect 3318 1348 3322 1352
rect 3342 1368 3346 1372
rect 3350 1348 3354 1352
rect 3342 1338 3346 1342
rect 3366 1338 3370 1342
rect 3358 1328 3362 1332
rect 3358 1308 3362 1312
rect 3398 1488 3402 1492
rect 3502 1658 3506 1662
rect 3510 1658 3514 1662
rect 3526 1648 3530 1652
rect 3654 1778 3658 1782
rect 3662 1778 3666 1782
rect 3542 1748 3546 1752
rect 3550 1748 3554 1752
rect 3566 1748 3570 1752
rect 3630 1748 3634 1752
rect 3590 1738 3594 1742
rect 3574 1708 3578 1712
rect 3542 1678 3546 1682
rect 3566 1678 3570 1682
rect 3598 1678 3602 1682
rect 3630 1698 3634 1702
rect 3638 1698 3642 1702
rect 3590 1668 3594 1672
rect 3574 1658 3578 1662
rect 3534 1638 3538 1642
rect 3502 1628 3506 1632
rect 3494 1618 3498 1622
rect 3494 1598 3498 1602
rect 3478 1578 3482 1582
rect 3470 1548 3474 1552
rect 3430 1518 3434 1522
rect 3470 1518 3474 1522
rect 3454 1478 3458 1482
rect 3446 1428 3450 1432
rect 3406 1418 3410 1422
rect 3410 1403 3414 1407
rect 3417 1403 3421 1407
rect 3398 1388 3402 1392
rect 3390 1358 3394 1362
rect 3622 1598 3626 1602
rect 3670 1768 3674 1772
rect 3678 1758 3682 1762
rect 3694 1748 3698 1752
rect 3678 1738 3682 1742
rect 3694 1738 3698 1742
rect 3686 1728 3690 1732
rect 3670 1698 3674 1702
rect 3646 1678 3650 1682
rect 3678 1678 3682 1682
rect 3670 1668 3674 1672
rect 3694 1668 3698 1672
rect 3702 1668 3706 1672
rect 3646 1658 3650 1662
rect 3662 1658 3666 1662
rect 3678 1658 3682 1662
rect 3694 1648 3698 1652
rect 3646 1628 3650 1632
rect 3670 1628 3674 1632
rect 3718 1758 3722 1762
rect 3766 1878 3770 1882
rect 3750 1858 3754 1862
rect 3742 1838 3746 1842
rect 3758 1838 3762 1842
rect 3742 1798 3746 1802
rect 3742 1768 3746 1772
rect 3734 1748 3738 1752
rect 3822 1838 3826 1842
rect 3774 1788 3778 1792
rect 3766 1758 3770 1762
rect 3758 1748 3762 1752
rect 3726 1688 3730 1692
rect 3766 1718 3770 1722
rect 3750 1708 3754 1712
rect 3718 1658 3722 1662
rect 3718 1648 3722 1652
rect 3726 1648 3730 1652
rect 3734 1638 3738 1642
rect 3750 1658 3754 1662
rect 3758 1648 3762 1652
rect 3742 1628 3746 1632
rect 3758 1628 3762 1632
rect 3710 1618 3714 1622
rect 3702 1598 3706 1602
rect 3542 1588 3546 1592
rect 3638 1588 3642 1592
rect 3502 1578 3506 1582
rect 3646 1578 3650 1582
rect 3494 1558 3498 1562
rect 3494 1548 3498 1552
rect 3486 1528 3490 1532
rect 3494 1498 3498 1502
rect 3494 1478 3498 1482
rect 3406 1348 3410 1352
rect 3446 1348 3450 1352
rect 3414 1328 3418 1332
rect 3406 1318 3410 1322
rect 3382 1298 3386 1302
rect 3350 1288 3354 1292
rect 3358 1288 3362 1292
rect 3342 1278 3346 1282
rect 3246 1268 3250 1272
rect 3270 1268 3274 1272
rect 3278 1268 3282 1272
rect 3318 1268 3322 1272
rect 3246 1258 3250 1262
rect 3142 1248 3146 1252
rect 3126 1168 3130 1172
rect 3038 1148 3042 1152
rect 3118 1148 3122 1152
rect 2998 1138 3002 1142
rect 3030 1138 3034 1142
rect 3062 1138 3066 1142
rect 2990 1128 2994 1132
rect 3006 1128 3010 1132
rect 3038 1128 3042 1132
rect 3062 1128 3066 1132
rect 3006 1118 3010 1122
rect 3030 1118 3034 1122
rect 3022 1108 3026 1112
rect 3078 1078 3082 1082
rect 2974 1068 2978 1072
rect 2958 1058 2962 1062
rect 3062 1058 3066 1062
rect 3078 1058 3082 1062
rect 2998 1048 3002 1052
rect 3014 1048 3018 1052
rect 2934 1038 2938 1042
rect 3022 1028 3026 1032
rect 3030 1028 3034 1032
rect 2918 1018 2922 1022
rect 2934 1018 2938 1022
rect 3014 1018 3018 1022
rect 2950 998 2954 1002
rect 2990 998 2994 1002
rect 2886 968 2890 972
rect 2958 968 2962 972
rect 3014 968 3018 972
rect 2910 958 2914 962
rect 2942 958 2946 962
rect 2878 948 2882 952
rect 2926 948 2930 952
rect 2982 948 2986 952
rect 2990 948 2994 952
rect 3006 948 3010 952
rect 2862 938 2866 942
rect 2830 928 2834 932
rect 2854 928 2858 932
rect 2814 918 2818 922
rect 2870 908 2874 912
rect 2830 898 2834 902
rect 2926 928 2930 932
rect 2906 903 2910 907
rect 2913 903 2917 907
rect 2846 878 2850 882
rect 2886 878 2890 882
rect 2918 878 2922 882
rect 2998 938 3002 942
rect 2958 908 2962 912
rect 2958 878 2962 882
rect 2990 918 2994 922
rect 2982 878 2986 882
rect 2838 868 2842 872
rect 2870 868 2874 872
rect 2902 868 2906 872
rect 2934 868 2938 872
rect 2966 868 2970 872
rect 2766 858 2770 862
rect 2782 858 2786 862
rect 2814 858 2818 862
rect 2766 838 2770 842
rect 2806 838 2810 842
rect 2758 818 2762 822
rect 2702 798 2706 802
rect 2702 768 2706 772
rect 2774 798 2778 802
rect 2694 748 2698 752
rect 2726 748 2730 752
rect 2758 748 2762 752
rect 2622 738 2626 742
rect 2734 738 2738 742
rect 2750 738 2754 742
rect 2798 768 2802 772
rect 2854 838 2858 842
rect 2894 838 2898 842
rect 2934 838 2938 842
rect 2846 788 2850 792
rect 2886 798 2890 802
rect 2862 778 2866 782
rect 2838 768 2842 772
rect 2854 768 2858 772
rect 2798 738 2802 742
rect 2670 728 2674 732
rect 2726 728 2730 732
rect 2774 728 2778 732
rect 2534 688 2538 692
rect 2526 668 2530 672
rect 2486 638 2490 642
rect 2510 638 2514 642
rect 2446 588 2450 592
rect 2446 558 2450 562
rect 2350 538 2354 542
rect 2390 498 2394 502
rect 2326 488 2330 492
rect 2318 478 2322 482
rect 2334 478 2338 482
rect 2366 478 2370 482
rect 2310 458 2314 462
rect 2342 458 2346 462
rect 2358 458 2362 462
rect 2374 458 2378 462
rect 2310 428 2314 432
rect 2342 398 2346 402
rect 2318 358 2322 362
rect 2342 348 2346 352
rect 2302 338 2306 342
rect 2342 338 2346 342
rect 2382 438 2386 442
rect 2374 408 2378 412
rect 2386 403 2390 407
rect 2393 403 2397 407
rect 2366 378 2370 382
rect 2374 378 2378 382
rect 2398 358 2402 362
rect 2366 348 2370 352
rect 2342 328 2346 332
rect 2262 318 2266 322
rect 2286 308 2290 312
rect 2302 288 2306 292
rect 2222 238 2226 242
rect 2270 238 2274 242
rect 2230 208 2234 212
rect 2182 188 2186 192
rect 2166 158 2170 162
rect 2134 148 2138 152
rect 2150 148 2154 152
rect 2158 148 2162 152
rect 2190 148 2194 152
rect 2126 138 2130 142
rect 2182 138 2186 142
rect 1918 128 1922 132
rect 2126 128 2130 132
rect 2006 108 2010 112
rect 1998 98 2002 102
rect 2094 88 2098 92
rect 2078 78 2082 82
rect 2038 68 2042 72
rect 2182 68 2186 72
rect 1966 58 1970 62
rect 2134 58 2138 62
rect 2238 158 2242 162
rect 2206 148 2210 152
rect 2270 198 2274 202
rect 2278 168 2282 172
rect 2278 148 2282 152
rect 2230 138 2234 142
rect 2246 138 2250 142
rect 2278 118 2282 122
rect 2206 108 2210 112
rect 2230 108 2234 112
rect 2214 88 2218 92
rect 2214 68 2218 72
rect 2294 108 2298 112
rect 2310 218 2314 222
rect 2382 328 2386 332
rect 2358 278 2362 282
rect 2350 208 2354 212
rect 2462 548 2466 552
rect 2454 498 2458 502
rect 2454 488 2458 492
rect 2414 478 2418 482
rect 2494 608 2498 612
rect 2470 488 2474 492
rect 2478 478 2482 482
rect 2486 478 2490 482
rect 2662 698 2666 702
rect 2726 698 2730 702
rect 2750 698 2754 702
rect 2734 688 2738 692
rect 2638 678 2642 682
rect 2686 678 2690 682
rect 2814 728 2818 732
rect 2814 708 2818 712
rect 2934 788 2938 792
rect 2910 768 2914 772
rect 2886 758 2890 762
rect 2878 748 2882 752
rect 2918 748 2922 752
rect 2830 738 2834 742
rect 2854 738 2858 742
rect 2862 738 2866 742
rect 2934 738 2938 742
rect 2990 858 2994 862
rect 2966 838 2970 842
rect 2950 808 2954 812
rect 3054 1018 3058 1022
rect 3038 978 3042 982
rect 3054 978 3058 982
rect 3030 928 3034 932
rect 3022 918 3026 922
rect 3078 978 3082 982
rect 3078 968 3082 972
rect 3134 1158 3138 1162
rect 3126 1118 3130 1122
rect 3102 1108 3106 1112
rect 3118 1108 3122 1112
rect 3094 1088 3098 1092
rect 3118 1088 3122 1092
rect 3166 1198 3170 1202
rect 3158 1158 3162 1162
rect 3158 1138 3162 1142
rect 3166 1138 3170 1142
rect 3142 1078 3146 1082
rect 3150 1068 3154 1072
rect 3102 1058 3106 1062
rect 3094 1048 3098 1052
rect 3110 1048 3114 1052
rect 3142 1048 3146 1052
rect 3102 1038 3106 1042
rect 3134 1038 3138 1042
rect 3150 968 3154 972
rect 3054 948 3058 952
rect 3086 948 3090 952
rect 3118 948 3122 952
rect 3134 948 3138 952
rect 3142 948 3146 952
rect 3070 938 3074 942
rect 3046 888 3050 892
rect 3030 868 3034 872
rect 3014 858 3018 862
rect 2950 778 2954 782
rect 2974 778 2978 782
rect 2934 728 2938 732
rect 2838 708 2842 712
rect 2846 698 2850 702
rect 2758 678 2762 682
rect 2838 678 2842 682
rect 2710 668 2714 672
rect 2774 668 2778 672
rect 2622 608 2626 612
rect 2582 598 2586 602
rect 2518 588 2522 592
rect 2726 598 2730 602
rect 2686 558 2690 562
rect 2718 558 2722 562
rect 2510 548 2514 552
rect 2622 548 2626 552
rect 2702 548 2706 552
rect 2718 548 2722 552
rect 2526 538 2530 542
rect 2558 518 2562 522
rect 2606 518 2610 522
rect 2622 518 2626 522
rect 2742 658 2746 662
rect 2790 658 2794 662
rect 2906 703 2910 707
rect 2913 703 2917 707
rect 2894 698 2898 702
rect 2854 688 2858 692
rect 2878 688 2882 692
rect 2894 688 2898 692
rect 2910 688 2914 692
rect 2886 668 2890 672
rect 2846 658 2850 662
rect 2958 768 2962 772
rect 2974 768 2978 772
rect 2958 738 2962 742
rect 3006 788 3010 792
rect 3086 918 3090 922
rect 3118 928 3122 932
rect 3134 928 3138 932
rect 3102 898 3106 902
rect 3126 888 3130 892
rect 3094 878 3098 882
rect 3102 868 3106 872
rect 3142 868 3146 872
rect 3110 858 3114 862
rect 3070 848 3074 852
rect 3054 838 3058 842
rect 3070 838 3074 842
rect 3086 838 3090 842
rect 3046 808 3050 812
rect 3022 768 3026 772
rect 3030 768 3034 772
rect 3014 748 3018 752
rect 2998 738 3002 742
rect 3022 738 3026 742
rect 2966 728 2970 732
rect 2982 728 2986 732
rect 3014 728 3018 732
rect 2990 698 2994 702
rect 2926 678 2930 682
rect 2974 658 2978 662
rect 2998 678 3002 682
rect 3054 738 3058 742
rect 3062 738 3066 742
rect 3038 708 3042 712
rect 3118 838 3122 842
rect 3102 818 3106 822
rect 3094 778 3098 782
rect 3078 768 3082 772
rect 3142 828 3146 832
rect 3166 1118 3170 1122
rect 3206 1238 3210 1242
rect 3190 1218 3194 1222
rect 3182 1198 3186 1202
rect 3222 1198 3226 1202
rect 3214 1188 3218 1192
rect 3270 1178 3274 1182
rect 3286 1248 3290 1252
rect 3302 1248 3306 1252
rect 3334 1228 3338 1232
rect 3182 1168 3186 1172
rect 3278 1168 3282 1172
rect 3374 1258 3378 1262
rect 3398 1308 3402 1312
rect 3414 1308 3418 1312
rect 3454 1308 3458 1312
rect 3422 1278 3426 1282
rect 3526 1568 3530 1572
rect 3542 1568 3546 1572
rect 3574 1568 3578 1572
rect 3622 1568 3626 1572
rect 3518 1548 3522 1552
rect 3534 1558 3538 1562
rect 3526 1538 3530 1542
rect 3558 1558 3562 1562
rect 3582 1558 3586 1562
rect 3614 1548 3618 1552
rect 3606 1538 3610 1542
rect 3638 1538 3642 1542
rect 3614 1528 3618 1532
rect 3550 1518 3554 1522
rect 3534 1478 3538 1482
rect 3574 1508 3578 1512
rect 3582 1498 3586 1502
rect 3558 1468 3562 1472
rect 3526 1458 3530 1462
rect 3502 1448 3506 1452
rect 3622 1518 3626 1522
rect 3638 1518 3642 1522
rect 3630 1498 3634 1502
rect 3590 1488 3594 1492
rect 3614 1478 3618 1482
rect 3590 1468 3594 1472
rect 3550 1448 3554 1452
rect 3558 1448 3562 1452
rect 3734 1568 3738 1572
rect 3654 1558 3658 1562
rect 3678 1548 3682 1552
rect 3670 1498 3674 1502
rect 3726 1558 3730 1562
rect 3710 1528 3714 1532
rect 3702 1488 3706 1492
rect 3654 1478 3658 1482
rect 3678 1478 3682 1482
rect 3686 1478 3690 1482
rect 3646 1468 3650 1472
rect 3662 1468 3666 1472
rect 3662 1448 3666 1452
rect 3622 1438 3626 1442
rect 3646 1428 3650 1432
rect 3566 1378 3570 1382
rect 3558 1368 3562 1372
rect 3550 1358 3554 1362
rect 3502 1348 3506 1352
rect 3526 1338 3530 1342
rect 3542 1338 3546 1342
rect 3574 1348 3578 1352
rect 3606 1348 3610 1352
rect 3622 1348 3626 1352
rect 3654 1348 3658 1352
rect 3566 1338 3570 1342
rect 3598 1338 3602 1342
rect 3614 1338 3618 1342
rect 3654 1338 3658 1342
rect 3478 1328 3482 1332
rect 3486 1318 3490 1322
rect 3510 1318 3514 1322
rect 3526 1318 3530 1322
rect 3478 1288 3482 1292
rect 3406 1268 3410 1272
rect 3414 1268 3418 1272
rect 3478 1268 3482 1272
rect 3390 1248 3394 1252
rect 3446 1248 3450 1252
rect 3422 1218 3426 1222
rect 3366 1178 3370 1182
rect 3410 1203 3414 1207
rect 3417 1203 3421 1207
rect 3534 1308 3538 1312
rect 3550 1308 3554 1312
rect 3542 1288 3546 1292
rect 3582 1328 3586 1332
rect 3622 1328 3626 1332
rect 3582 1308 3586 1312
rect 3670 1308 3674 1312
rect 3646 1298 3650 1302
rect 3582 1288 3586 1292
rect 3598 1288 3602 1292
rect 3494 1268 3498 1272
rect 3502 1238 3506 1242
rect 3486 1208 3490 1212
rect 3534 1248 3538 1252
rect 3510 1188 3514 1192
rect 3550 1188 3554 1192
rect 3374 1168 3378 1172
rect 3206 1158 3210 1162
rect 3254 1158 3258 1162
rect 3326 1158 3330 1162
rect 3342 1158 3346 1162
rect 3470 1158 3474 1162
rect 3222 1148 3226 1152
rect 3190 1138 3194 1142
rect 3182 1108 3186 1112
rect 3190 1078 3194 1082
rect 3174 998 3178 1002
rect 3182 968 3186 972
rect 3238 1138 3242 1142
rect 3366 1148 3370 1152
rect 3454 1148 3458 1152
rect 3326 1138 3330 1142
rect 3230 1128 3234 1132
rect 3246 1128 3250 1132
rect 3278 1128 3282 1132
rect 3246 1118 3250 1122
rect 3302 1118 3306 1122
rect 3230 1098 3234 1102
rect 3334 1088 3338 1092
rect 3246 1078 3250 1082
rect 3350 1138 3354 1142
rect 3382 1128 3386 1132
rect 3222 1068 3226 1072
rect 3286 1068 3290 1072
rect 3342 1068 3346 1072
rect 3358 1068 3362 1072
rect 3206 1058 3210 1062
rect 3238 1058 3242 1062
rect 3230 1048 3234 1052
rect 3310 1058 3314 1062
rect 3286 1048 3290 1052
rect 3446 1138 3450 1142
rect 3462 1138 3466 1142
rect 3478 1138 3482 1142
rect 3494 1178 3498 1182
rect 3550 1168 3554 1172
rect 3422 1128 3426 1132
rect 3454 1128 3458 1132
rect 3470 1128 3474 1132
rect 3486 1128 3490 1132
rect 3430 1118 3434 1122
rect 3438 1108 3442 1112
rect 3494 1118 3498 1122
rect 3526 1148 3530 1152
rect 3510 1128 3514 1132
rect 3518 1108 3522 1112
rect 3462 1088 3466 1092
rect 3470 1078 3474 1082
rect 3430 1068 3434 1072
rect 3374 1058 3378 1062
rect 3406 1058 3410 1062
rect 3438 1058 3442 1062
rect 3350 1048 3354 1052
rect 3214 1028 3218 1032
rect 3262 1028 3266 1032
rect 3294 1028 3298 1032
rect 3342 1028 3346 1032
rect 3198 1018 3202 1022
rect 3198 958 3202 962
rect 3174 938 3178 942
rect 3166 928 3170 932
rect 3158 898 3162 902
rect 3166 888 3170 892
rect 3166 858 3170 862
rect 3174 848 3178 852
rect 3318 1008 3322 1012
rect 3310 988 3314 992
rect 3230 958 3234 962
rect 3262 948 3266 952
rect 3294 948 3298 952
rect 3310 948 3314 952
rect 3206 878 3210 882
rect 3198 868 3202 872
rect 3230 898 3234 902
rect 3278 938 3282 942
rect 3302 938 3306 942
rect 3246 928 3250 932
rect 3262 928 3266 932
rect 3286 928 3290 932
rect 3294 908 3298 912
rect 3302 888 3306 892
rect 3262 868 3266 872
rect 3214 858 3218 862
rect 3246 858 3250 862
rect 3206 848 3210 852
rect 3254 848 3258 852
rect 3158 838 3162 842
rect 3182 818 3186 822
rect 3150 808 3154 812
rect 3142 768 3146 772
rect 3110 758 3114 762
rect 3134 758 3138 762
rect 3086 738 3090 742
rect 3118 728 3122 732
rect 3126 718 3130 722
rect 3134 718 3138 722
rect 3078 688 3082 692
rect 3110 688 3114 692
rect 3102 668 3106 672
rect 3118 668 3122 672
rect 3006 658 3010 662
rect 3046 658 3050 662
rect 2758 638 2762 642
rect 2782 638 2786 642
rect 2830 638 2834 642
rect 2886 638 2890 642
rect 2910 638 2914 642
rect 2974 638 2978 642
rect 2742 598 2746 602
rect 2766 568 2770 572
rect 2798 568 2802 572
rect 2942 608 2946 612
rect 2878 598 2882 602
rect 2766 558 2770 562
rect 2870 558 2874 562
rect 2742 548 2746 552
rect 2886 568 2890 572
rect 2958 568 2962 572
rect 2774 548 2778 552
rect 2870 548 2874 552
rect 2886 548 2890 552
rect 2918 548 2922 552
rect 2942 548 2946 552
rect 2694 538 2698 542
rect 2734 538 2738 542
rect 2798 538 2802 542
rect 2814 538 2818 542
rect 2966 558 2970 562
rect 2974 548 2978 552
rect 2638 478 2642 482
rect 2654 478 2658 482
rect 2662 478 2666 482
rect 2494 468 2498 472
rect 2590 468 2594 472
rect 2430 458 2434 462
rect 2446 458 2450 462
rect 2454 458 2458 462
rect 2438 428 2442 432
rect 2422 398 2426 402
rect 2502 458 2506 462
rect 2494 438 2498 442
rect 2534 438 2538 442
rect 2574 438 2578 442
rect 2590 438 2594 442
rect 2502 428 2506 432
rect 2414 388 2418 392
rect 2446 388 2450 392
rect 2462 388 2466 392
rect 2414 358 2418 362
rect 2462 358 2466 362
rect 2494 358 2498 362
rect 2526 418 2530 422
rect 2518 368 2522 372
rect 2438 348 2442 352
rect 2422 338 2426 342
rect 2406 328 2410 332
rect 2422 328 2426 332
rect 2470 348 2474 352
rect 2502 348 2506 352
rect 2510 338 2514 342
rect 2390 298 2394 302
rect 2438 288 2442 292
rect 2630 458 2634 462
rect 2630 438 2634 442
rect 2614 428 2618 432
rect 2582 408 2586 412
rect 2558 398 2562 402
rect 2590 398 2594 402
rect 2606 398 2610 402
rect 2582 388 2586 392
rect 2646 468 2650 472
rect 2646 438 2650 442
rect 2750 528 2754 532
rect 2718 478 2722 482
rect 2822 528 2826 532
rect 2838 528 2842 532
rect 2822 518 2826 522
rect 2790 498 2794 502
rect 2814 498 2818 502
rect 2830 498 2834 502
rect 2710 468 2714 472
rect 2742 468 2746 472
rect 2774 468 2778 472
rect 2750 458 2754 462
rect 2758 448 2762 452
rect 2686 438 2690 442
rect 2742 398 2746 402
rect 2742 388 2746 392
rect 2694 368 2698 372
rect 2766 368 2770 372
rect 2702 358 2706 362
rect 2734 358 2738 362
rect 2766 358 2770 362
rect 2670 348 2674 352
rect 2694 348 2698 352
rect 2718 348 2722 352
rect 2542 308 2546 312
rect 2558 308 2562 312
rect 2582 308 2586 312
rect 2550 298 2554 302
rect 2566 298 2570 302
rect 2478 248 2482 252
rect 2386 203 2390 207
rect 2393 203 2397 207
rect 2430 188 2434 192
rect 2470 188 2474 192
rect 2502 248 2506 252
rect 2534 228 2538 232
rect 2622 298 2626 302
rect 2590 278 2594 282
rect 2574 268 2578 272
rect 2590 268 2594 272
rect 2870 528 2874 532
rect 2918 528 2922 532
rect 2894 518 2898 522
rect 2822 488 2826 492
rect 2846 488 2850 492
rect 2870 478 2874 482
rect 2846 468 2850 472
rect 2798 448 2802 452
rect 2870 458 2874 462
rect 2838 448 2842 452
rect 2846 448 2850 452
rect 2870 448 2874 452
rect 2822 438 2826 442
rect 2814 418 2818 422
rect 2782 388 2786 392
rect 2750 348 2754 352
rect 2774 348 2778 352
rect 2702 338 2706 342
rect 2710 338 2714 342
rect 2758 338 2762 342
rect 2678 298 2682 302
rect 2686 298 2690 302
rect 2702 298 2706 302
rect 2614 258 2618 262
rect 2590 248 2594 252
rect 2558 208 2562 212
rect 2574 198 2578 202
rect 2358 158 2362 162
rect 2398 158 2402 162
rect 2486 158 2490 162
rect 2518 158 2522 162
rect 2342 148 2346 152
rect 2558 138 2562 142
rect 2630 238 2634 242
rect 2646 228 2650 232
rect 2630 188 2634 192
rect 2662 238 2666 242
rect 2654 188 2658 192
rect 2774 218 2778 222
rect 2718 178 2722 182
rect 2742 178 2746 182
rect 2710 158 2714 162
rect 2726 148 2730 152
rect 2694 138 2698 142
rect 2734 138 2738 142
rect 2678 128 2682 132
rect 2646 108 2650 112
rect 2294 98 2298 102
rect 2302 98 2306 102
rect 2374 98 2378 102
rect 2606 98 2610 102
rect 2582 88 2586 92
rect 2758 78 2762 82
rect 2294 68 2298 72
rect 2494 68 2498 72
rect 2670 68 2674 72
rect 2798 368 2802 372
rect 2830 368 2834 372
rect 2822 358 2826 362
rect 2790 348 2794 352
rect 2862 358 2866 362
rect 2906 503 2910 507
rect 2913 503 2917 507
rect 2910 468 2914 472
rect 2942 478 2946 482
rect 2990 638 2994 642
rect 2990 558 2994 562
rect 3014 638 3018 642
rect 3062 638 3066 642
rect 3014 558 3018 562
rect 3030 558 3034 562
rect 3054 558 3058 562
rect 3014 548 3018 552
rect 2998 538 3002 542
rect 3070 538 3074 542
rect 3022 508 3026 512
rect 3062 528 3066 532
rect 3110 628 3114 632
rect 3110 578 3114 582
rect 3118 568 3122 572
rect 3094 558 3098 562
rect 3142 638 3146 642
rect 3142 558 3146 562
rect 3126 548 3130 552
rect 3086 538 3090 542
rect 3078 518 3082 522
rect 3038 498 3042 502
rect 3070 498 3074 502
rect 3046 478 3050 482
rect 2974 468 2978 472
rect 2894 438 2898 442
rect 2894 398 2898 402
rect 2854 348 2858 352
rect 2878 348 2882 352
rect 2926 458 2930 462
rect 2950 458 2954 462
rect 2974 458 2978 462
rect 3022 458 3026 462
rect 2942 448 2946 452
rect 2990 448 2994 452
rect 2918 368 2922 372
rect 2966 438 2970 442
rect 3014 428 3018 432
rect 2974 388 2978 392
rect 3046 448 3050 452
rect 3038 388 3042 392
rect 2982 378 2986 382
rect 2974 368 2978 372
rect 2934 358 2938 362
rect 3014 358 3018 362
rect 2918 348 2922 352
rect 2822 328 2826 332
rect 2886 328 2890 332
rect 2854 318 2858 322
rect 2878 318 2882 322
rect 2906 303 2910 307
rect 2913 303 2917 307
rect 2870 298 2874 302
rect 2862 278 2866 282
rect 2846 268 2850 272
rect 2790 258 2794 262
rect 2838 258 2842 262
rect 2838 238 2842 242
rect 2846 238 2850 242
rect 2830 218 2834 222
rect 2830 148 2834 152
rect 2958 328 2962 332
rect 2950 308 2954 312
rect 2902 248 2906 252
rect 2886 238 2890 242
rect 2878 218 2882 222
rect 2894 218 2898 222
rect 2870 208 2874 212
rect 2846 138 2850 142
rect 2798 128 2802 132
rect 2822 128 2826 132
rect 2846 118 2850 122
rect 2854 98 2858 102
rect 2854 88 2858 92
rect 2886 148 2890 152
rect 2886 78 2890 82
rect 2934 278 2938 282
rect 2990 298 2994 302
rect 2982 268 2986 272
rect 2934 258 2938 262
rect 2910 198 2914 202
rect 2942 248 2946 252
rect 3014 278 3018 282
rect 3022 268 3026 272
rect 3014 258 3018 262
rect 3014 248 3018 252
rect 2974 228 2978 232
rect 2982 228 2986 232
rect 2974 178 2978 182
rect 2958 168 2962 172
rect 2942 158 2946 162
rect 2966 148 2970 152
rect 3038 288 3042 292
rect 3142 528 3146 532
rect 3134 488 3138 492
rect 3182 768 3186 772
rect 3174 758 3178 762
rect 3214 838 3218 842
rect 3238 838 3242 842
rect 3230 788 3234 792
rect 3230 768 3234 772
rect 3262 758 3266 762
rect 3390 1048 3394 1052
rect 3454 1048 3458 1052
rect 3406 1038 3410 1042
rect 3398 1028 3402 1032
rect 3366 968 3370 972
rect 3334 948 3338 952
rect 3358 948 3362 952
rect 3318 878 3322 882
rect 3326 868 3330 872
rect 3350 938 3354 942
rect 3366 938 3370 942
rect 3382 958 3386 962
rect 3502 1068 3506 1072
rect 3494 1048 3498 1052
rect 3502 1038 3506 1042
rect 3486 1018 3490 1022
rect 3410 1003 3414 1007
rect 3417 1003 3421 1007
rect 3422 978 3426 982
rect 3494 978 3498 982
rect 3398 948 3402 952
rect 3510 988 3514 992
rect 3470 968 3474 972
rect 3502 968 3506 972
rect 3446 928 3450 932
rect 3470 908 3474 912
rect 3406 888 3410 892
rect 3374 878 3378 882
rect 3510 958 3514 962
rect 3486 948 3490 952
rect 3502 948 3506 952
rect 3542 1098 3546 1102
rect 3582 1268 3586 1272
rect 3606 1268 3610 1272
rect 3566 1258 3570 1262
rect 3582 1258 3586 1262
rect 3678 1298 3682 1302
rect 3678 1288 3682 1292
rect 3638 1258 3642 1262
rect 3662 1258 3666 1262
rect 3678 1258 3682 1262
rect 3574 1238 3578 1242
rect 3566 1168 3570 1172
rect 3558 1148 3562 1152
rect 3614 1238 3618 1242
rect 3638 1228 3642 1232
rect 3622 1218 3626 1222
rect 3630 1208 3634 1212
rect 3582 1158 3586 1162
rect 3550 1078 3554 1082
rect 3566 1078 3570 1082
rect 3534 1068 3538 1072
rect 3558 1068 3562 1072
rect 3550 1058 3554 1062
rect 3606 1178 3610 1182
rect 3614 1158 3618 1162
rect 3614 1138 3618 1142
rect 3630 1128 3634 1132
rect 3598 1108 3602 1112
rect 3598 1088 3602 1092
rect 3590 1078 3594 1082
rect 3526 998 3530 1002
rect 3606 1068 3610 1072
rect 3614 1068 3618 1072
rect 3590 1038 3594 1042
rect 3614 1038 3618 1042
rect 3622 1038 3626 1042
rect 3582 978 3586 982
rect 3614 1028 3618 1032
rect 3630 1018 3634 1022
rect 3606 978 3610 982
rect 3590 968 3594 972
rect 3518 938 3522 942
rect 3526 938 3530 942
rect 3510 918 3514 922
rect 3526 898 3530 902
rect 3518 888 3522 892
rect 3342 868 3346 872
rect 3406 868 3410 872
rect 3454 868 3458 872
rect 3510 868 3514 872
rect 3334 858 3338 862
rect 3350 858 3354 862
rect 3462 858 3466 862
rect 3478 858 3482 862
rect 3342 848 3346 852
rect 3358 848 3362 852
rect 3382 848 3386 852
rect 3318 838 3322 842
rect 3350 838 3354 842
rect 3278 748 3282 752
rect 3190 738 3194 742
rect 3262 738 3266 742
rect 3206 728 3210 732
rect 3230 728 3234 732
rect 3246 728 3250 732
rect 3158 718 3162 722
rect 3174 718 3178 722
rect 3254 708 3258 712
rect 3214 698 3218 702
rect 3158 678 3162 682
rect 3214 678 3218 682
rect 3262 688 3266 692
rect 3158 658 3162 662
rect 3198 658 3202 662
rect 3238 658 3242 662
rect 3222 648 3226 652
rect 3158 608 3162 612
rect 3190 608 3194 612
rect 3182 598 3186 602
rect 3174 568 3178 572
rect 3182 558 3186 562
rect 3158 548 3162 552
rect 3166 548 3170 552
rect 3286 678 3290 682
rect 3334 748 3338 752
rect 3454 848 3458 852
rect 3470 848 3474 852
rect 3398 838 3402 842
rect 3446 838 3450 842
rect 3410 803 3414 807
rect 3417 803 3421 807
rect 3438 788 3442 792
rect 3462 768 3466 772
rect 3382 758 3386 762
rect 3518 848 3522 852
rect 3486 838 3490 842
rect 3486 758 3490 762
rect 3390 748 3394 752
rect 3478 748 3482 752
rect 3310 738 3314 742
rect 3318 728 3322 732
rect 3334 728 3338 732
rect 3302 718 3306 722
rect 3310 688 3314 692
rect 3310 658 3314 662
rect 3270 638 3274 642
rect 3254 578 3258 582
rect 3214 568 3218 572
rect 3238 568 3242 572
rect 3214 538 3218 542
rect 3222 538 3226 542
rect 3254 558 3258 562
rect 3190 528 3194 532
rect 3230 498 3234 502
rect 3238 478 3242 482
rect 3358 738 3362 742
rect 3398 738 3402 742
rect 3470 738 3474 742
rect 3374 728 3378 732
rect 3382 718 3386 722
rect 3422 728 3426 732
rect 3446 728 3450 732
rect 3462 718 3466 722
rect 3518 818 3522 822
rect 3550 958 3554 962
rect 3558 928 3562 932
rect 3622 958 3626 962
rect 3574 918 3578 922
rect 3590 918 3594 922
rect 3582 908 3586 912
rect 3558 888 3562 892
rect 3582 878 3586 882
rect 3566 858 3570 862
rect 3558 848 3562 852
rect 3574 848 3578 852
rect 3590 838 3594 842
rect 3598 828 3602 832
rect 3646 1158 3650 1162
rect 3646 1128 3650 1132
rect 3646 1058 3650 1062
rect 3646 1038 3650 1042
rect 3670 1228 3674 1232
rect 3662 1038 3666 1042
rect 3654 1018 3658 1022
rect 3702 1468 3706 1472
rect 3718 1458 3722 1462
rect 3718 1438 3722 1442
rect 3694 1428 3698 1432
rect 3710 1418 3714 1422
rect 3702 1378 3706 1382
rect 3742 1548 3746 1552
rect 3758 1458 3762 1462
rect 3758 1448 3762 1452
rect 3750 1438 3754 1442
rect 3726 1418 3730 1422
rect 3742 1418 3746 1422
rect 3734 1408 3738 1412
rect 3726 1378 3730 1382
rect 3758 1398 3762 1402
rect 3742 1368 3746 1372
rect 3774 1638 3778 1642
rect 3766 1388 3770 1392
rect 3774 1368 3778 1372
rect 3766 1358 3770 1362
rect 3710 1348 3714 1352
rect 3766 1348 3770 1352
rect 3694 1338 3698 1342
rect 3750 1328 3754 1332
rect 3694 1318 3698 1322
rect 3726 1298 3730 1302
rect 3702 1278 3706 1282
rect 3718 1278 3722 1282
rect 3758 1288 3762 1292
rect 3742 1278 3746 1282
rect 3726 1268 3730 1272
rect 3726 1258 3730 1262
rect 3758 1258 3762 1262
rect 3734 1248 3738 1252
rect 3750 1248 3754 1252
rect 3694 1238 3698 1242
rect 3822 1218 3826 1222
rect 3758 1198 3762 1202
rect 3726 1178 3730 1182
rect 3750 1168 3754 1172
rect 3742 1148 3746 1152
rect 3726 1138 3730 1142
rect 3742 1138 3746 1142
rect 3686 1098 3690 1102
rect 3686 1088 3690 1092
rect 3702 1078 3706 1082
rect 3734 1078 3738 1082
rect 3678 1068 3682 1072
rect 3710 1058 3714 1062
rect 3694 998 3698 1002
rect 3662 988 3666 992
rect 3646 968 3650 972
rect 3670 958 3674 962
rect 3686 958 3690 962
rect 3622 928 3626 932
rect 3638 878 3642 882
rect 3638 868 3642 872
rect 3670 928 3674 932
rect 3718 1028 3722 1032
rect 3726 938 3730 942
rect 3718 928 3722 932
rect 3686 908 3690 912
rect 3694 908 3698 912
rect 3710 908 3714 912
rect 3630 848 3634 852
rect 3622 828 3626 832
rect 3638 808 3642 812
rect 3622 788 3626 792
rect 3542 778 3546 782
rect 3502 768 3506 772
rect 3510 748 3514 752
rect 3502 738 3506 742
rect 3510 698 3514 702
rect 3478 688 3482 692
rect 3486 688 3490 692
rect 3358 678 3362 682
rect 3422 678 3426 682
rect 3334 658 3338 662
rect 3374 658 3378 662
rect 3326 648 3330 652
rect 3286 638 3290 642
rect 3342 628 3346 632
rect 3286 598 3290 602
rect 3302 558 3306 562
rect 3278 538 3282 542
rect 3270 528 3274 532
rect 3398 658 3402 662
rect 3438 658 3442 662
rect 3390 608 3394 612
rect 3410 603 3414 607
rect 3417 603 3421 607
rect 3342 598 3346 602
rect 3334 568 3338 572
rect 3382 578 3386 582
rect 3350 548 3354 552
rect 3326 538 3330 542
rect 3342 538 3346 542
rect 3262 518 3266 522
rect 3294 518 3298 522
rect 3358 518 3362 522
rect 3350 498 3354 502
rect 3302 478 3306 482
rect 3326 478 3330 482
rect 3190 468 3194 472
rect 3262 468 3266 472
rect 3094 458 3098 462
rect 3078 388 3082 392
rect 3102 388 3106 392
rect 3150 368 3154 372
rect 3094 358 3098 362
rect 3150 358 3154 362
rect 3166 358 3170 362
rect 3078 338 3082 342
rect 3110 318 3114 322
rect 3110 308 3114 312
rect 3102 248 3106 252
rect 3158 338 3162 342
rect 3230 458 3234 462
rect 3222 398 3226 402
rect 3214 368 3218 372
rect 3198 338 3202 342
rect 3230 338 3234 342
rect 3134 328 3138 332
rect 3174 328 3178 332
rect 3182 328 3186 332
rect 3150 298 3154 302
rect 3206 278 3210 282
rect 3150 268 3154 272
rect 3190 268 3194 272
rect 3190 258 3194 262
rect 3142 248 3146 252
rect 3126 228 3130 232
rect 3054 208 3058 212
rect 3030 198 3034 202
rect 3062 198 3066 202
rect 3006 188 3010 192
rect 3070 188 3074 192
rect 3086 208 3090 212
rect 3006 158 3010 162
rect 3038 158 3042 162
rect 3078 158 3082 162
rect 2990 148 2994 152
rect 3006 148 3010 152
rect 2926 138 2930 142
rect 2998 138 3002 142
rect 3022 138 3026 142
rect 3046 138 3050 142
rect 3006 128 3010 132
rect 2906 103 2910 107
rect 2913 103 2917 107
rect 3022 118 3026 122
rect 3102 198 3106 202
rect 3094 118 3098 122
rect 3094 88 3098 92
rect 3510 678 3514 682
rect 3630 778 3634 782
rect 3550 758 3554 762
rect 3582 758 3586 762
rect 3606 758 3610 762
rect 3542 688 3546 692
rect 3574 718 3578 722
rect 3566 708 3570 712
rect 3574 698 3578 702
rect 3534 668 3538 672
rect 3478 648 3482 652
rect 3454 628 3458 632
rect 3462 618 3466 622
rect 3454 608 3458 612
rect 3438 548 3442 552
rect 3614 728 3618 732
rect 3606 708 3610 712
rect 3614 708 3618 712
rect 3606 688 3610 692
rect 3598 668 3602 672
rect 3558 658 3562 662
rect 3566 658 3570 662
rect 3518 648 3522 652
rect 3510 608 3514 612
rect 3574 648 3578 652
rect 3582 648 3586 652
rect 3598 618 3602 622
rect 3654 878 3658 882
rect 3662 868 3666 872
rect 3686 868 3690 872
rect 3702 868 3706 872
rect 3670 858 3674 862
rect 3646 788 3650 792
rect 3702 838 3706 842
rect 3718 868 3722 872
rect 3758 958 3762 962
rect 3774 1118 3778 1122
rect 3774 1068 3778 1072
rect 3774 948 3778 952
rect 3750 928 3754 932
rect 3742 858 3746 862
rect 3702 828 3706 832
rect 3710 828 3714 832
rect 3686 798 3690 802
rect 3686 788 3690 792
rect 3654 778 3658 782
rect 3670 778 3674 782
rect 3686 768 3690 772
rect 3654 748 3658 752
rect 3670 748 3674 752
rect 3686 748 3690 752
rect 3686 728 3690 732
rect 3646 718 3650 722
rect 3630 698 3634 702
rect 3566 568 3570 572
rect 3598 568 3602 572
rect 3470 558 3474 562
rect 3614 558 3618 562
rect 3494 548 3498 552
rect 3518 548 3522 552
rect 3534 548 3538 552
rect 3558 548 3562 552
rect 3574 548 3578 552
rect 3606 548 3610 552
rect 3518 538 3522 542
rect 3422 528 3426 532
rect 3446 528 3450 532
rect 3478 528 3482 532
rect 3510 528 3514 532
rect 3406 518 3410 522
rect 3582 538 3586 542
rect 3598 538 3602 542
rect 3542 528 3546 532
rect 3534 518 3538 522
rect 3494 508 3498 512
rect 3398 498 3402 502
rect 3574 518 3578 522
rect 3382 488 3386 492
rect 3534 488 3538 492
rect 3446 478 3450 482
rect 3534 478 3538 482
rect 3366 468 3370 472
rect 3374 468 3378 472
rect 3462 468 3466 472
rect 3270 458 3274 462
rect 3286 448 3290 452
rect 3270 438 3274 442
rect 3254 408 3258 412
rect 3302 378 3306 382
rect 3278 348 3282 352
rect 3254 308 3258 312
rect 3302 338 3306 342
rect 3278 318 3282 322
rect 3294 318 3298 322
rect 3350 438 3354 442
rect 3334 408 3338 412
rect 3326 358 3330 362
rect 3286 308 3290 312
rect 3310 308 3314 312
rect 3270 298 3274 302
rect 3278 298 3282 302
rect 3270 278 3274 282
rect 3334 338 3338 342
rect 3318 288 3322 292
rect 3350 358 3354 362
rect 3390 448 3394 452
rect 3382 418 3386 422
rect 3446 438 3450 442
rect 3410 403 3414 407
rect 3417 403 3421 407
rect 3510 418 3514 422
rect 3486 368 3490 372
rect 3462 358 3466 362
rect 3358 348 3362 352
rect 3438 348 3442 352
rect 3478 348 3482 352
rect 3382 338 3386 342
rect 3430 338 3434 342
rect 3470 338 3474 342
rect 3350 328 3354 332
rect 3374 328 3378 332
rect 3414 328 3418 332
rect 3462 308 3466 312
rect 3406 298 3410 302
rect 3446 288 3450 292
rect 3326 278 3330 282
rect 3246 268 3250 272
rect 3334 268 3338 272
rect 3278 258 3282 262
rect 3318 258 3322 262
rect 3302 238 3306 242
rect 3302 228 3306 232
rect 3278 218 3282 222
rect 3326 248 3330 252
rect 3310 198 3314 202
rect 3238 178 3242 182
rect 3158 148 3162 152
rect 3142 138 3146 142
rect 3126 108 3130 112
rect 3110 98 3114 102
rect 3142 88 3146 92
rect 2990 78 2994 82
rect 3142 78 3146 82
rect 3222 138 3226 142
rect 3286 138 3290 142
rect 3302 138 3306 142
rect 3230 128 3234 132
rect 3246 78 3250 82
rect 3046 68 3050 72
rect 3190 68 3194 72
rect 3310 118 3314 122
rect 3638 628 3642 632
rect 3662 658 3666 662
rect 3686 648 3690 652
rect 3678 628 3682 632
rect 3654 608 3658 612
rect 3734 828 3738 832
rect 3726 788 3730 792
rect 3726 778 3730 782
rect 3750 768 3754 772
rect 3766 758 3770 762
rect 3710 738 3714 742
rect 3710 718 3714 722
rect 3718 708 3722 712
rect 3710 678 3714 682
rect 3726 668 3730 672
rect 3726 648 3730 652
rect 3702 638 3706 642
rect 3694 618 3698 622
rect 3686 608 3690 612
rect 3646 558 3650 562
rect 3646 538 3650 542
rect 3630 508 3634 512
rect 3582 488 3586 492
rect 3678 558 3682 562
rect 3670 498 3674 502
rect 3670 488 3674 492
rect 3598 468 3602 472
rect 3614 468 3618 472
rect 3646 468 3650 472
rect 3590 458 3594 462
rect 3558 418 3562 422
rect 3518 358 3522 362
rect 3502 348 3506 352
rect 3582 438 3586 442
rect 3574 338 3578 342
rect 3518 318 3522 322
rect 3502 278 3506 282
rect 3502 268 3506 272
rect 3454 208 3458 212
rect 3410 203 3414 207
rect 3417 203 3421 207
rect 3406 188 3410 192
rect 3422 148 3426 152
rect 3366 138 3370 142
rect 3406 138 3410 142
rect 3398 98 3402 102
rect 3334 68 3338 72
rect 3358 68 3362 72
rect 3390 68 3394 72
rect 2222 58 2226 62
rect 2510 58 2514 62
rect 2566 58 2570 62
rect 2630 58 2634 62
rect 2686 58 2690 62
rect 2742 58 2746 62
rect 2782 58 2786 62
rect 2830 58 2834 62
rect 2846 58 2850 62
rect 2910 58 2914 62
rect 2950 58 2954 62
rect 3126 58 3130 62
rect 3366 58 3370 62
rect 1998 28 2002 32
rect 1926 8 1930 12
rect 2406 48 2410 52
rect 3494 248 3498 252
rect 3534 218 3538 222
rect 3534 208 3538 212
rect 3542 178 3546 182
rect 3446 88 3450 92
rect 3430 78 3434 82
rect 3486 78 3490 82
rect 3470 68 3474 72
rect 3558 168 3562 172
rect 3566 168 3570 172
rect 3550 148 3554 152
rect 3622 448 3626 452
rect 3654 448 3658 452
rect 3614 438 3618 442
rect 3638 438 3642 442
rect 3606 428 3610 432
rect 3606 408 3610 412
rect 3598 318 3602 322
rect 3590 288 3594 292
rect 3590 188 3594 192
rect 3598 158 3602 162
rect 3574 118 3578 122
rect 3630 428 3634 432
rect 3702 598 3706 602
rect 3694 548 3698 552
rect 3710 548 3714 552
rect 3718 538 3722 542
rect 3710 518 3714 522
rect 3718 518 3722 522
rect 3694 508 3698 512
rect 3702 508 3706 512
rect 3702 488 3706 492
rect 3686 468 3690 472
rect 3718 508 3722 512
rect 3758 748 3762 752
rect 3750 688 3754 692
rect 3758 678 3762 682
rect 3742 658 3746 662
rect 3750 648 3754 652
rect 3766 648 3770 652
rect 3750 638 3754 642
rect 3734 578 3738 582
rect 3766 568 3770 572
rect 3742 528 3746 532
rect 3742 498 3746 502
rect 3734 488 3738 492
rect 3710 468 3714 472
rect 3734 468 3738 472
rect 3694 458 3698 462
rect 3726 458 3730 462
rect 3718 428 3722 432
rect 3646 368 3650 372
rect 3614 358 3618 362
rect 3630 358 3634 362
rect 3654 358 3658 362
rect 3662 358 3666 362
rect 3758 348 3762 352
rect 3622 338 3626 342
rect 3638 328 3642 332
rect 3622 318 3626 322
rect 3614 258 3618 262
rect 3606 108 3610 112
rect 3598 88 3602 92
rect 3622 148 3626 152
rect 3646 318 3650 322
rect 3646 298 3650 302
rect 3630 88 3634 92
rect 3550 68 3554 72
rect 3590 68 3594 72
rect 3662 338 3666 342
rect 3702 338 3706 342
rect 3758 318 3762 322
rect 3694 288 3698 292
rect 3710 278 3714 282
rect 3710 248 3714 252
rect 3718 218 3722 222
rect 3766 228 3770 232
rect 3758 208 3762 212
rect 3742 198 3746 202
rect 3718 168 3722 172
rect 3662 158 3666 162
rect 3718 158 3722 162
rect 3678 148 3682 152
rect 3670 138 3674 142
rect 3662 128 3666 132
rect 3702 128 3706 132
rect 3694 108 3698 112
rect 3686 88 3690 92
rect 3718 98 3722 102
rect 3734 88 3738 92
rect 3718 78 3722 82
rect 3678 68 3682 72
rect 3694 68 3698 72
rect 3478 58 3482 62
rect 3526 58 3530 62
rect 3614 58 3618 62
rect 3654 58 3658 62
rect 3686 58 3690 62
rect 3710 58 3714 62
rect 3758 78 3762 82
rect 3358 48 3362 52
rect 3646 48 3650 52
rect 3726 48 3730 52
rect 3334 38 3338 42
rect 3374 38 3378 42
rect 3390 38 3394 42
rect 3454 38 3458 42
rect 3590 38 3594 42
rect 3750 38 3754 42
rect 3342 28 3346 32
rect 2094 8 2098 12
rect 2494 8 2498 12
rect 2386 3 2390 7
rect 2393 3 2397 7
rect 3410 3 3414 7
rect 3417 3 3421 7
<< metal3 >>
rect 344 3603 346 3607
rect 350 3603 353 3607
rect 358 3603 360 3607
rect 1360 3603 1362 3607
rect 1366 3603 1369 3607
rect 1374 3603 1376 3607
rect 2384 3603 2386 3607
rect 2390 3603 2393 3607
rect 2398 3603 2400 3607
rect 3408 3603 3410 3607
rect 3414 3603 3417 3607
rect 3422 3603 3424 3607
rect 426 3598 430 3601
rect 890 3598 894 3601
rect 1466 3598 1478 3601
rect 1506 3598 1510 3601
rect 1962 3598 1974 3601
rect 1070 3592 1073 3598
rect 1334 3592 1337 3598
rect 1574 3592 1577 3598
rect 1606 3592 1609 3598
rect 1758 3592 1761 3598
rect 1902 3592 1905 3598
rect 2230 3592 2233 3598
rect 2406 3592 2409 3598
rect 1274 3588 1278 3591
rect 1502 3588 1510 3591
rect 1514 3588 1526 3591
rect 1794 3588 1798 3591
rect 2074 3588 2078 3591
rect 2434 3588 2902 3591
rect 2906 3588 2942 3591
rect 2946 3588 2974 3591
rect 3118 3588 3262 3591
rect 3266 3588 3334 3591
rect 3118 3582 3121 3588
rect 1386 3578 1398 3581
rect 1590 3578 2766 3581
rect 3342 3581 3345 3588
rect 3242 3578 3345 3581
rect 1590 3572 1593 3578
rect 1082 3568 1590 3571
rect 2066 3568 2070 3571
rect 2266 3568 2454 3571
rect 3198 3571 3201 3578
rect 2954 3568 3201 3571
rect 3322 3568 3342 3571
rect 3458 3568 3478 3571
rect 3482 3568 3534 3571
rect 3682 3568 3686 3571
rect 1866 3558 2022 3561
rect 2026 3558 2126 3561
rect 2130 3558 2366 3561
rect 2410 3558 2446 3561
rect 2478 3561 2481 3568
rect 2474 3558 2481 3561
rect 2754 3558 2910 3561
rect 3178 3558 3230 3561
rect 3234 3558 3438 3561
rect 3442 3558 3462 3561
rect 3466 3558 3502 3561
rect 3662 3552 3665 3558
rect 322 3548 374 3551
rect 522 3548 606 3551
rect 730 3548 734 3551
rect 1154 3548 1206 3551
rect 1394 3548 1470 3551
rect 1994 3548 2190 3551
rect 2514 3548 2854 3551
rect 2898 3548 2926 3551
rect 3186 3548 3222 3551
rect 3250 3548 3278 3551
rect 3338 3548 3350 3551
rect 3354 3548 3374 3551
rect 3378 3548 3390 3551
rect 3434 3548 3454 3551
rect 3466 3548 3470 3551
rect 3538 3548 3566 3551
rect 3610 3548 3614 3551
rect 1662 3542 1665 3548
rect 34 3538 62 3541
rect 66 3538 86 3541
rect 90 3538 102 3541
rect 106 3538 174 3541
rect 662 3538 670 3541
rect 1122 3538 1238 3541
rect 1354 3538 1486 3541
rect 1574 3538 1582 3541
rect 2002 3538 2006 3541
rect 2162 3538 2166 3541
rect 2362 3538 2382 3541
rect 2422 3541 2425 3548
rect 3150 3542 3153 3548
rect 2402 3538 2470 3541
rect 2634 3538 2702 3541
rect 2810 3538 2974 3541
rect 3210 3538 3214 3541
rect 3286 3541 3289 3548
rect 3326 3542 3329 3548
rect 3286 3538 3310 3541
rect 3482 3538 3550 3541
rect 3658 3538 3662 3541
rect 3738 3538 3745 3541
rect 662 3532 665 3538
rect 902 3532 905 3538
rect 1062 3532 1065 3538
rect 1574 3532 1577 3538
rect 1798 3532 1801 3538
rect 242 3528 449 3531
rect 962 3528 966 3531
rect 1634 3528 1750 3531
rect 1814 3531 1817 3538
rect 1814 3528 1854 3531
rect 2014 3531 2017 3538
rect 2278 3532 2281 3538
rect 2574 3532 2577 3538
rect 1986 3528 2166 3531
rect 2194 3528 2262 3531
rect 2490 3528 2494 3531
rect 2834 3528 3022 3531
rect 3154 3528 3254 3531
rect 3446 3531 3449 3538
rect 3742 3532 3745 3538
rect 3266 3528 3449 3531
rect 3650 3528 3710 3531
rect 3730 3528 3734 3531
rect 446 3522 449 3528
rect 1302 3522 1305 3528
rect 1974 3522 1977 3528
rect 290 3518 294 3521
rect 450 3518 702 3521
rect 706 3518 886 3521
rect 1234 3518 1286 3521
rect 2178 3518 2430 3521
rect 2858 3518 2926 3521
rect 2946 3518 3038 3521
rect 3154 3518 3294 3521
rect 3298 3518 3334 3521
rect 3354 3518 3382 3521
rect 3386 3518 3478 3521
rect 3510 3521 3513 3528
rect 3598 3522 3601 3528
rect 3510 3518 3558 3521
rect 426 3508 430 3511
rect 874 3508 1078 3511
rect 1146 3508 1166 3511
rect 1306 3508 1398 3511
rect 1906 3508 1982 3511
rect 2234 3508 2238 3511
rect 2250 3508 2270 3511
rect 2282 3508 2438 3511
rect 2442 3508 2462 3511
rect 2530 3508 2670 3511
rect 2674 3508 2870 3511
rect 3082 3508 3158 3511
rect 3194 3508 3254 3511
rect 3266 3508 3294 3511
rect 3298 3508 3566 3511
rect 848 3503 850 3507
rect 854 3503 857 3507
rect 862 3503 864 3507
rect 1286 3502 1289 3508
rect 1880 3503 1882 3507
rect 1886 3503 1889 3507
rect 1894 3503 1896 3507
rect 2904 3503 2906 3507
rect 2910 3503 2913 3507
rect 2918 3503 2920 3507
rect 1334 3498 1438 3501
rect 1954 3498 1966 3501
rect 2042 3498 2438 3501
rect 2442 3498 2590 3501
rect 2930 3498 2998 3501
rect 3002 3498 3158 3501
rect 3162 3498 3278 3501
rect 3282 3498 3310 3501
rect 3314 3498 3542 3501
rect 3546 3498 3590 3501
rect 3650 3498 3758 3501
rect 538 3488 646 3491
rect 650 3488 689 3491
rect 1270 3488 1278 3491
rect 1334 3491 1337 3498
rect 1282 3488 1337 3491
rect 1346 3488 1374 3491
rect 1442 3488 1990 3491
rect 1994 3488 2038 3491
rect 2098 3488 2142 3491
rect 2186 3488 2254 3491
rect 2274 3488 2566 3491
rect 3042 3488 3118 3491
rect 3218 3488 3518 3491
rect 3586 3488 3598 3491
rect 3610 3488 3694 3491
rect 170 3478 678 3481
rect 686 3481 689 3488
rect 686 3478 1742 3481
rect 1882 3478 2886 3481
rect 2890 3478 2894 3481
rect 2902 3481 2905 3488
rect 2902 3478 3118 3481
rect 3122 3478 3302 3481
rect 3306 3478 3462 3481
rect 3510 3478 3518 3481
rect 3522 3478 3566 3481
rect 3586 3478 3606 3481
rect 3722 3478 3729 3481
rect 318 3472 321 3478
rect 1614 3472 1617 3478
rect 334 3468 702 3471
rect 1226 3468 1246 3471
rect 1250 3468 1270 3471
rect 1274 3468 1302 3471
rect 1814 3471 1817 3478
rect 3726 3472 3729 3478
rect 3742 3472 3745 3478
rect 1814 3468 1902 3471
rect 2006 3468 2022 3471
rect 2202 3468 2238 3471
rect 2306 3468 2537 3471
rect 2546 3468 2574 3471
rect 2578 3468 2582 3471
rect 2802 3468 2809 3471
rect 2866 3468 2878 3471
rect 2938 3468 3358 3471
rect 3362 3468 3438 3471
rect 3482 3468 3510 3471
rect 3514 3468 3582 3471
rect 3634 3468 3670 3471
rect 6 3462 9 3468
rect 334 3462 337 3468
rect 894 3462 897 3468
rect 1422 3462 1425 3468
rect 2006 3462 2009 3468
rect 2534 3462 2537 3468
rect 610 3458 630 3461
rect 1218 3458 1262 3461
rect 1266 3458 1286 3461
rect 1290 3458 1310 3461
rect 1482 3458 1526 3461
rect 1530 3458 1542 3461
rect 2130 3458 2190 3461
rect 2226 3458 2254 3461
rect 2266 3458 2270 3461
rect 2554 3458 2558 3461
rect 2578 3458 2798 3461
rect 2806 3461 2809 3468
rect 2806 3458 3009 3461
rect 3018 3458 3070 3461
rect 3114 3458 3382 3461
rect 3394 3458 3430 3461
rect 3442 3458 3526 3461
rect 3554 3458 3566 3461
rect 3626 3458 3686 3461
rect 198 3452 201 3458
rect 3006 3452 3009 3458
rect 3702 3452 3705 3458
rect -26 3451 -22 3452
rect -26 3448 6 3451
rect 442 3448 646 3451
rect 662 3448 1222 3451
rect 1754 3448 2150 3451
rect 2194 3448 2214 3451
rect 2530 3448 2542 3451
rect 2562 3448 2758 3451
rect 2762 3448 2886 3451
rect 2962 3448 2966 3451
rect 3018 3448 3134 3451
rect 3138 3448 3190 3451
rect 3210 3448 3214 3451
rect 3234 3448 3270 3451
rect 3290 3448 3502 3451
rect 3642 3448 3678 3451
rect 662 3441 665 3448
rect 562 3438 665 3441
rect 994 3438 1262 3441
rect 1866 3438 2046 3441
rect 2166 3441 2169 3448
rect 3590 3442 3593 3448
rect 3774 3442 3777 3448
rect 2166 3438 2334 3441
rect 2338 3438 2814 3441
rect 2818 3438 2846 3441
rect 2850 3438 2870 3441
rect 2882 3438 2974 3441
rect 2986 3438 3030 3441
rect 3034 3438 3142 3441
rect 3242 3438 3254 3441
rect 3266 3438 3494 3441
rect 3530 3438 3534 3441
rect 3538 3438 3558 3441
rect 3618 3438 3630 3441
rect 3658 3438 3662 3441
rect 138 3428 582 3431
rect 586 3428 870 3431
rect 1058 3428 1081 3431
rect 1162 3428 1190 3431
rect 1194 3428 1318 3431
rect 1518 3431 1521 3438
rect 1518 3428 2558 3431
rect 2982 3431 2985 3438
rect 2754 3428 2985 3431
rect 3142 3431 3145 3438
rect 3670 3432 3673 3438
rect 3142 3428 3462 3431
rect 3466 3428 3518 3431
rect 3522 3428 3542 3431
rect 3546 3428 3654 3431
rect 86 3421 89 3428
rect 86 3418 942 3421
rect 1066 3418 1070 3421
rect 1078 3421 1081 3428
rect 1078 3418 1270 3421
rect 1610 3418 1614 3421
rect 1858 3418 1870 3421
rect 1874 3418 2086 3421
rect 2226 3418 2302 3421
rect 2306 3418 2414 3421
rect 2530 3418 2662 3421
rect 2786 3418 2934 3421
rect 2938 3418 3062 3421
rect 3066 3418 3166 3421
rect 3178 3418 3246 3421
rect 3258 3418 3262 3421
rect 3274 3418 3278 3421
rect 3290 3418 3414 3421
rect 3542 3418 3550 3421
rect 3554 3418 3606 3421
rect 3702 3421 3705 3428
rect 3674 3418 3705 3421
rect 178 3408 294 3411
rect 554 3408 598 3411
rect 674 3408 734 3411
rect 1058 3408 1318 3411
rect 1386 3408 2182 3411
rect 2186 3408 2374 3411
rect 2458 3408 2622 3411
rect 2834 3408 2990 3411
rect 3226 3408 3286 3411
rect 3298 3408 3302 3411
rect 3458 3408 3542 3411
rect 3578 3408 3750 3411
rect 344 3403 346 3407
rect 350 3403 353 3407
rect 358 3403 360 3407
rect 1360 3403 1362 3407
rect 1366 3403 1369 3407
rect 1374 3403 1376 3407
rect 2384 3403 2386 3407
rect 2390 3403 2393 3407
rect 2398 3403 2400 3407
rect 3408 3403 3410 3407
rect 3414 3403 3417 3407
rect 3422 3403 3424 3407
rect 26 3398 326 3401
rect 458 3398 558 3401
rect 658 3398 1246 3401
rect 1250 3398 1342 3401
rect 1578 3398 1582 3401
rect 1722 3398 1750 3401
rect 1802 3398 1910 3401
rect 2954 3398 3374 3401
rect 3506 3398 3630 3401
rect 3698 3398 3734 3401
rect 186 3388 238 3391
rect 242 3388 286 3391
rect 290 3388 318 3391
rect 362 3388 382 3391
rect 386 3388 409 3391
rect 978 3388 1086 3391
rect 1306 3388 1406 3391
rect 1626 3388 1798 3391
rect 1802 3388 2006 3391
rect 2090 3388 2278 3391
rect 2282 3388 2294 3391
rect 2646 3391 2649 3398
rect 2646 3388 2958 3391
rect 2986 3388 3198 3391
rect 3250 3388 3326 3391
rect 3346 3388 3430 3391
rect 3434 3388 3478 3391
rect 3490 3388 3598 3391
rect 3602 3388 3678 3391
rect 406 3382 409 3388
rect 890 3378 998 3381
rect 1306 3378 1478 3381
rect 1622 3381 1625 3388
rect 1482 3378 1625 3381
rect 1746 3378 2526 3381
rect 2874 3378 2950 3381
rect 2954 3378 3006 3381
rect 3010 3378 3014 3381
rect 3026 3378 3182 3381
rect 3194 3378 3270 3381
rect 3282 3378 3366 3381
rect 3378 3378 3614 3381
rect 3618 3378 3670 3381
rect 3722 3378 3726 3381
rect -26 3371 -22 3372
rect 6 3371 9 3378
rect -26 3368 9 3371
rect 250 3368 454 3371
rect 882 3368 1230 3371
rect 1322 3368 1590 3371
rect 1602 3368 1622 3371
rect 1658 3368 2358 3371
rect 2362 3368 2550 3371
rect 2778 3368 3094 3371
rect 3098 3368 3190 3371
rect 3194 3368 3222 3371
rect 3250 3368 3254 3371
rect 3298 3368 3302 3371
rect 3322 3368 3342 3371
rect 3354 3368 3582 3371
rect 3586 3368 3598 3371
rect 3602 3368 3630 3371
rect 3730 3368 3774 3371
rect 1310 3362 1313 3368
rect -26 3358 30 3361
rect 354 3358 870 3361
rect 954 3358 1262 3361
rect 1266 3358 1297 3361
rect 1378 3358 1982 3361
rect 1986 3358 1993 3361
rect 2002 3358 2390 3361
rect 2394 3358 2406 3361
rect 2890 3358 2894 3361
rect 2970 3358 2998 3361
rect 3002 3358 3022 3361
rect 3058 3358 3206 3361
rect 3234 3358 3270 3361
rect 3346 3358 3374 3361
rect 3418 3358 3422 3361
rect 3426 3358 3510 3361
rect 3522 3358 3558 3361
rect 3562 3358 3590 3361
rect 3594 3358 3622 3361
rect 3698 3358 3718 3361
rect -26 3352 -23 3358
rect 1294 3352 1297 3358
rect -26 3348 -22 3352
rect 26 3348 246 3351
rect 322 3348 366 3351
rect 426 3348 878 3351
rect 946 3348 1046 3351
rect 1114 3348 1126 3351
rect 1242 3348 1262 3351
rect 1314 3348 1358 3351
rect 1378 3348 1558 3351
rect 1754 3348 1798 3351
rect 1930 3348 2174 3351
rect 2178 3348 2318 3351
rect 2370 3348 2486 3351
rect 2878 3351 2881 3358
rect 3126 3352 3129 3358
rect 2682 3348 2881 3351
rect 2930 3348 3014 3351
rect 3170 3348 3278 3351
rect 3290 3348 3310 3351
rect 3370 3348 3382 3351
rect 3490 3348 3518 3351
rect 3530 3348 3550 3351
rect 3610 3348 3646 3351
rect 3650 3348 3686 3351
rect 58 3338 70 3341
rect 314 3338 398 3341
rect 610 3338 774 3341
rect 786 3338 830 3341
rect 834 3338 982 3341
rect 994 3338 1022 3341
rect 1042 3338 1110 3341
rect 1274 3338 1326 3341
rect 1354 3338 1358 3341
rect 1426 3338 1497 3341
rect 1602 3338 1774 3341
rect 1850 3338 1857 3341
rect 1494 3332 1497 3338
rect 1854 3332 1857 3338
rect 2170 3338 2782 3341
rect 2890 3338 2902 3341
rect 2970 3338 2998 3341
rect 3114 3338 3134 3341
rect 3138 3338 3246 3341
rect 3334 3341 3337 3348
rect 3334 3338 3406 3341
rect 3410 3338 3454 3341
rect 3682 3338 3686 3341
rect 3714 3338 3718 3341
rect 3722 3338 3750 3341
rect 2110 3332 2113 3338
rect 66 3328 254 3331
rect 274 3328 281 3331
rect 394 3328 446 3331
rect 450 3328 614 3331
rect 682 3328 785 3331
rect 850 3328 902 3331
rect 954 3328 974 3331
rect 1194 3328 1318 3331
rect 1610 3328 1678 3331
rect 2194 3328 2198 3331
rect 2306 3328 2310 3331
rect 2594 3328 2606 3331
rect 2610 3328 2678 3331
rect 2898 3328 2926 3331
rect 2978 3328 3174 3331
rect 3294 3331 3297 3338
rect 3274 3328 3350 3331
rect 3354 3328 3382 3331
rect 3498 3328 3526 3331
rect 3674 3328 3718 3331
rect 3746 3328 3758 3331
rect 178 3318 262 3321
rect 278 3321 281 3328
rect 782 3322 785 3328
rect 266 3318 273 3321
rect 278 3318 414 3321
rect 506 3318 518 3321
rect 538 3318 662 3321
rect 786 3318 1070 3321
rect 1074 3318 1182 3321
rect 1194 3318 1382 3321
rect 1394 3318 1398 3321
rect 1482 3318 1590 3321
rect 1786 3318 1974 3321
rect 1978 3318 2126 3321
rect 2226 3318 2246 3321
rect 2306 3318 2358 3321
rect 2362 3318 2382 3321
rect 2426 3318 2449 3321
rect 2802 3318 2953 3321
rect 3010 3318 3046 3321
rect 3066 3318 3102 3321
rect 3206 3321 3209 3328
rect 3206 3318 3270 3321
rect 3282 3318 3318 3321
rect 3374 3318 3382 3321
rect 3386 3318 3438 3321
rect 3442 3318 3462 3321
rect 3638 3321 3641 3328
rect 3626 3318 3641 3321
rect 3662 3321 3665 3328
rect 3662 3318 3758 3321
rect 2446 3312 2449 3318
rect 2950 3312 2953 3318
rect 178 3308 206 3311
rect 282 3308 550 3311
rect 634 3308 694 3311
rect 706 3308 774 3311
rect 890 3308 926 3311
rect 1290 3308 1350 3311
rect 1354 3308 1510 3311
rect 1514 3308 1862 3311
rect 2026 3308 2318 3311
rect 2498 3308 2542 3311
rect 2674 3308 2870 3311
rect 2954 3308 2982 3311
rect 2986 3308 3030 3311
rect 3090 3308 3174 3311
rect 3266 3308 3278 3311
rect 3402 3308 3678 3311
rect 3682 3308 3734 3311
rect 848 3303 850 3307
rect 854 3303 857 3307
rect 862 3303 864 3307
rect 1880 3303 1882 3307
rect 1886 3303 1889 3307
rect 1894 3303 1896 3307
rect 2014 3302 2017 3308
rect 2904 3303 2906 3307
rect 2910 3303 2913 3307
rect 2918 3303 2920 3307
rect 226 3298 230 3301
rect 234 3298 286 3301
rect 290 3298 318 3301
rect 322 3298 366 3301
rect 378 3298 470 3301
rect 474 3298 622 3301
rect 626 3298 646 3301
rect 690 3298 766 3301
rect 874 3298 982 3301
rect 986 3298 1022 3301
rect 1090 3298 1134 3301
rect 1330 3298 1689 3301
rect 1698 3298 1758 3301
rect 2102 3298 2694 3301
rect 2930 3298 3014 3301
rect 3042 3298 3070 3301
rect 3250 3298 3334 3301
rect 3538 3298 3646 3301
rect 3650 3298 3662 3301
rect 3666 3298 3726 3301
rect 410 3288 518 3291
rect 1242 3288 1326 3291
rect 1338 3288 1382 3291
rect 1402 3288 1414 3291
rect 1418 3288 1462 3291
rect 1506 3288 1510 3291
rect 1686 3291 1689 3298
rect 1686 3288 1702 3291
rect 2102 3291 2105 3298
rect 1874 3288 2105 3291
rect 2898 3288 3038 3291
rect 3122 3288 3150 3291
rect 3154 3288 3230 3291
rect 3234 3288 3246 3291
rect 3346 3288 3478 3291
rect 3546 3288 3614 3291
rect 370 3278 478 3281
rect 954 3278 1206 3281
rect 1210 3278 1262 3281
rect 1410 3278 1486 3281
rect 1634 3278 1662 3281
rect 1666 3278 1686 3281
rect 1690 3278 1694 3281
rect 1790 3281 1793 3288
rect 1786 3278 1793 3281
rect 2182 3281 2185 3288
rect 2098 3278 2185 3281
rect 2298 3278 2342 3281
rect 2410 3278 2438 3281
rect 2506 3278 2518 3281
rect 2522 3278 2566 3281
rect 2782 3281 2785 3288
rect 2782 3278 2854 3281
rect 2874 3278 2918 3281
rect 2922 3278 3006 3281
rect 3018 3278 3038 3281
rect 3098 3278 3166 3281
rect 3178 3278 3182 3281
rect 3186 3278 3238 3281
rect 3250 3278 3342 3281
rect 3402 3278 3462 3281
rect 3522 3278 3550 3281
rect 3638 3281 3641 3288
rect 3638 3278 3686 3281
rect 3698 3278 3742 3281
rect 782 3272 785 3278
rect 942 3272 945 3278
rect 3766 3272 3769 3278
rect 290 3268 510 3271
rect 562 3268 606 3271
rect 690 3268 702 3271
rect 786 3268 806 3271
rect 946 3268 1110 3271
rect 1114 3268 1158 3271
rect 1266 3268 1310 3271
rect 1330 3268 1638 3271
rect 1658 3268 1678 3271
rect 1682 3268 1806 3271
rect 1810 3268 1902 3271
rect 2130 3268 2366 3271
rect 2370 3268 2510 3271
rect 2650 3268 2801 3271
rect 2906 3268 2926 3271
rect 2930 3268 2950 3271
rect 2970 3268 2974 3271
rect 3010 3268 3014 3271
rect 3018 3268 3062 3271
rect 3090 3268 3158 3271
rect 3226 3268 3278 3271
rect 3306 3268 3350 3271
rect 3354 3268 3550 3271
rect 3610 3268 3638 3271
rect 134 3262 137 3268
rect 450 3258 454 3261
rect 610 3258 622 3261
rect 678 3261 681 3268
rect 626 3258 681 3261
rect 714 3258 814 3261
rect 1018 3258 1038 3261
rect 1226 3258 1230 3261
rect 1234 3258 1286 3261
rect 1298 3258 1302 3261
rect 1338 3258 1398 3261
rect 2306 3258 2342 3261
rect 2394 3258 2414 3261
rect 2450 3258 2486 3261
rect 2546 3258 2550 3261
rect 2598 3261 2601 3268
rect 2578 3258 2601 3261
rect 2798 3262 2801 3268
rect 3174 3262 3177 3268
rect 2962 3258 2982 3261
rect 2986 3258 3014 3261
rect 3026 3258 3054 3261
rect 3102 3258 3126 3261
rect 3290 3258 3318 3261
rect 3322 3258 3358 3261
rect 3370 3258 3374 3261
rect 3378 3258 3398 3261
rect 3410 3258 3422 3261
rect 3490 3258 3510 3261
rect 3546 3258 3550 3261
rect 3554 3258 3574 3261
rect 3618 3258 3646 3261
rect 3698 3258 3718 3261
rect 1094 3252 1097 3258
rect 3102 3252 3105 3258
rect -26 3251 -22 3252
rect -26 3248 6 3251
rect 122 3248 134 3251
rect 138 3248 318 3251
rect 442 3248 510 3251
rect 514 3248 534 3251
rect 562 3248 566 3251
rect 594 3248 598 3251
rect 762 3248 766 3251
rect 1306 3248 1358 3251
rect 1410 3248 1446 3251
rect 1490 3248 1510 3251
rect 1542 3248 1870 3251
rect 1890 3248 1894 3251
rect 2286 3248 2310 3251
rect 2370 3248 2470 3251
rect 2474 3248 2590 3251
rect 2634 3248 2694 3251
rect 2890 3248 2918 3251
rect 2922 3248 3062 3251
rect 3154 3248 3182 3251
rect 3234 3248 3294 3251
rect 3330 3248 3390 3251
rect 3394 3248 3438 3251
rect 3530 3248 3542 3251
rect 3554 3248 3710 3251
rect 3766 3251 3769 3258
rect 3730 3248 3769 3251
rect 1262 3242 1265 3248
rect 114 3238 206 3241
rect 426 3238 478 3241
rect 530 3238 718 3241
rect 722 3238 742 3241
rect 1274 3238 1310 3241
rect 1398 3241 1401 3248
rect 1542 3242 1545 3248
rect 2286 3242 2289 3248
rect 3238 3242 3241 3248
rect 1314 3238 1401 3241
rect 1410 3238 1542 3241
rect 1554 3238 2166 3241
rect 2378 3238 2390 3241
rect 2482 3238 2494 3241
rect 3042 3238 3126 3241
rect 3162 3238 3182 3241
rect 3202 3238 3230 3241
rect 3506 3238 3534 3241
rect 3554 3238 3582 3241
rect 3594 3238 3718 3241
rect 1270 3232 1273 3238
rect 306 3228 721 3231
rect 1234 3228 1262 3231
rect 1290 3228 1334 3231
rect 1530 3228 1750 3231
rect 2194 3228 2270 3231
rect 2274 3228 2438 3231
rect 2442 3228 2510 3231
rect 2514 3228 2566 3231
rect 2726 3228 3718 3231
rect 3722 3228 3766 3231
rect 718 3222 721 3228
rect 210 3218 630 3221
rect 2726 3221 2729 3228
rect 1170 3218 2729 3221
rect 3082 3218 3206 3221
rect 3210 3218 3310 3221
rect 3314 3218 3374 3221
rect 3706 3218 3718 3221
rect 966 3212 969 3218
rect 458 3208 486 3211
rect 1402 3208 1454 3211
rect 1458 3208 1558 3211
rect 1770 3208 1798 3211
rect 1802 3208 2294 3211
rect 2298 3208 2310 3211
rect 3130 3208 3270 3211
rect 344 3203 346 3207
rect 350 3203 353 3207
rect 358 3203 360 3207
rect 1360 3203 1362 3207
rect 1366 3203 1369 3207
rect 1374 3203 1376 3207
rect 1710 3202 1713 3208
rect 2384 3203 2386 3207
rect 2390 3203 2393 3207
rect 2398 3203 2400 3207
rect 3408 3203 3410 3207
rect 3414 3203 3417 3207
rect 3422 3203 3424 3207
rect 682 3198 694 3201
rect 1306 3198 1342 3201
rect 1810 3198 1886 3201
rect 1930 3198 1934 3201
rect 2026 3198 2038 3201
rect 2066 3198 2102 3201
rect 2178 3198 2198 3201
rect 2298 3198 2310 3201
rect 2746 3198 2758 3201
rect 3266 3198 3366 3201
rect 322 3188 1174 3191
rect 1178 3188 1278 3191
rect 1322 3188 1726 3191
rect 1834 3188 1846 3191
rect 2338 3188 2502 3191
rect 3058 3188 3286 3191
rect 3594 3188 3678 3191
rect 578 3178 582 3181
rect 778 3178 830 3181
rect 834 3178 886 3181
rect 1354 3178 1526 3181
rect 1618 3178 2438 3181
rect 2442 3178 2622 3181
rect 2626 3178 2670 3181
rect 3282 3178 3350 3181
rect 3554 3178 3702 3181
rect 3158 3172 3161 3178
rect 754 3168 798 3171
rect 802 3168 878 3171
rect 918 3168 926 3171
rect 930 3168 974 3171
rect 1538 3168 1790 3171
rect 1814 3168 1929 3171
rect 1938 3168 1966 3171
rect 2002 3168 2110 3171
rect 2214 3168 2294 3171
rect 2362 3168 2390 3171
rect 2418 3168 2606 3171
rect 2610 3168 2630 3171
rect 2866 3168 2926 3171
rect 3262 3171 3265 3178
rect 3262 3168 3542 3171
rect 3570 3168 3686 3171
rect 3690 3168 3710 3171
rect 218 3158 726 3161
rect 746 3158 766 3161
rect 770 3158 798 3161
rect 802 3158 870 3161
rect 982 3161 985 3168
rect 882 3158 985 3161
rect 1002 3158 1006 3161
rect 1266 3158 1414 3161
rect 1418 3158 1430 3161
rect 1494 3161 1497 3168
rect 1798 3162 1801 3168
rect 1814 3162 1817 3168
rect 1494 3158 1518 3161
rect 1530 3158 1614 3161
rect 1646 3158 1686 3161
rect 1690 3158 1710 3161
rect 1874 3158 1902 3161
rect 1906 3158 1910 3161
rect 1926 3161 1929 3168
rect 2214 3162 2217 3168
rect 1926 3158 2062 3161
rect 2066 3158 2078 3161
rect 2090 3158 2150 3161
rect 2154 3158 2201 3161
rect 2226 3158 2230 3161
rect 2354 3158 2398 3161
rect 2514 3158 2526 3161
rect 2566 3158 2590 3161
rect 2926 3161 2929 3168
rect 2926 3158 3078 3161
rect 3138 3158 3142 3161
rect 3154 3158 3166 3161
rect 3178 3158 3206 3161
rect 3322 3158 3334 3161
rect 3354 3158 3382 3161
rect 3402 3158 3430 3161
rect 3506 3158 3526 3161
rect 3554 3158 3598 3161
rect 3626 3158 3630 3161
rect 3634 3158 3726 3161
rect 282 3148 294 3151
rect 298 3148 366 3151
rect 522 3148 526 3151
rect 706 3148 814 3151
rect 842 3148 918 3151
rect 922 3148 958 3151
rect 1010 3148 1014 3151
rect 1130 3148 1142 3151
rect 1146 3148 1206 3151
rect 1266 3148 1422 3151
rect 1458 3148 1486 3151
rect 1646 3151 1649 3158
rect 2158 3152 2161 3158
rect 2198 3152 2201 3158
rect 2566 3152 2569 3158
rect 1642 3148 1649 3151
rect 1658 3148 1838 3151
rect 1842 3148 1854 3151
rect 1962 3148 1974 3151
rect 1978 3148 1985 3151
rect 1994 3148 2022 3151
rect 2050 3148 2070 3151
rect 2226 3148 2254 3151
rect 2298 3148 2422 3151
rect 2426 3148 2454 3151
rect 2522 3148 2542 3151
rect 2586 3148 2638 3151
rect 3018 3148 3174 3151
rect 3182 3148 3286 3151
rect 3290 3148 3326 3151
rect 3358 3148 3438 3151
rect 3474 3148 3502 3151
rect 3570 3148 3574 3151
rect 3618 3148 3662 3151
rect -26 3141 -22 3142
rect -26 3138 6 3141
rect 10 3138 14 3141
rect 406 3141 409 3148
rect 406 3138 526 3141
rect 582 3141 585 3148
rect 974 3142 977 3148
rect 582 3138 718 3141
rect 730 3138 846 3141
rect 914 3138 934 3141
rect 938 3138 942 3141
rect 986 3138 1318 3141
rect 1418 3138 1462 3141
rect 1514 3138 1582 3141
rect 1586 3138 1694 3141
rect 1698 3138 1782 3141
rect 1898 3138 1926 3141
rect 1938 3138 2118 3141
rect 2178 3138 2214 3141
rect 2298 3138 2302 3141
rect 2318 3138 2438 3141
rect 2442 3138 2518 3141
rect 2602 3138 2606 3141
rect 3182 3141 3185 3148
rect 3358 3142 3361 3148
rect 3002 3138 3185 3141
rect 3194 3138 3257 3141
rect 3394 3138 3406 3141
rect 3450 3138 3478 3141
rect 3490 3138 3534 3141
rect 3610 3138 3654 3141
rect 2318 3132 2321 3138
rect 170 3128 502 3131
rect 714 3128 734 3131
rect 762 3128 766 3131
rect 778 3128 942 3131
rect 946 3128 1193 3131
rect 1202 3128 1406 3131
rect 1410 3128 1438 3131
rect 1482 3128 1630 3131
rect 1634 3128 1782 3131
rect 1786 3128 1798 3131
rect 1842 3128 1942 3131
rect 1946 3128 1966 3131
rect 2018 3128 2038 3131
rect 2114 3128 2126 3131
rect 2130 3128 2222 3131
rect 2242 3128 2246 3131
rect 2330 3128 2366 3131
rect 2466 3128 2470 3131
rect 2474 3128 2510 3131
rect 2566 3131 2569 3138
rect 2774 3132 2777 3138
rect 3254 3132 3257 3138
rect 2566 3128 2758 3131
rect 3034 3128 3094 3131
rect 3138 3128 3150 3131
rect 3306 3128 3342 3131
rect 3346 3128 3398 3131
rect 3442 3128 3518 3131
rect 3742 3131 3745 3138
rect 3658 3128 3745 3131
rect 230 3122 233 3128
rect 422 3122 425 3128
rect 598 3122 601 3128
rect 746 3118 758 3121
rect 826 3118 950 3121
rect 1190 3121 1193 3128
rect 1190 3118 1542 3121
rect 1738 3118 1742 3121
rect 1798 3121 1801 3128
rect 1798 3118 1942 3121
rect 1946 3118 1982 3121
rect 1994 3118 2022 3121
rect 2066 3118 2118 3121
rect 2234 3118 2454 3121
rect 2594 3118 2598 3121
rect 2682 3118 2934 3121
rect 2938 3118 2990 3121
rect 3158 3121 3161 3128
rect 3114 3118 3161 3121
rect 3218 3118 3262 3121
rect 3590 3121 3593 3128
rect 3590 3118 3678 3121
rect 3682 3118 3726 3121
rect 1614 3112 1617 3118
rect 1758 3112 1761 3118
rect 578 3108 782 3111
rect 1098 3108 1102 3111
rect 1474 3108 1542 3111
rect 1682 3108 1750 3111
rect 2054 3111 2057 3118
rect 1938 3108 2057 3111
rect 2122 3108 2222 3111
rect 2250 3108 2262 3111
rect 2266 3108 2310 3111
rect 2322 3108 2686 3111
rect 2690 3108 2702 3111
rect 3122 3108 3134 3111
rect 3202 3108 3214 3111
rect 848 3103 850 3107
rect 854 3103 857 3107
rect 862 3103 864 3107
rect 1880 3103 1882 3107
rect 1886 3103 1889 3107
rect 1894 3103 1896 3107
rect 2904 3103 2906 3107
rect 2910 3103 2913 3107
rect 2918 3103 2920 3107
rect 258 3098 310 3101
rect 314 3098 774 3101
rect 1090 3098 1246 3101
rect 1250 3098 1406 3101
rect 1698 3098 1710 3101
rect 1714 3098 1822 3101
rect 1986 3098 2118 3101
rect 2130 3098 2150 3101
rect 2250 3098 2254 3101
rect 2290 3098 2398 3101
rect 2538 3098 2590 3101
rect 2594 3098 2622 3101
rect 2634 3098 2662 3101
rect 3098 3098 3113 3101
rect 3122 3098 3230 3101
rect 3234 3098 3302 3101
rect 3306 3098 3374 3101
rect 1870 3092 1873 3098
rect 1354 3088 1526 3091
rect 1554 3088 1601 3091
rect 1618 3088 1678 3091
rect 2018 3088 2030 3091
rect 2034 3088 2278 3091
rect 2306 3088 2422 3091
rect 2490 3088 2806 3091
rect 2810 3088 2862 3091
rect 3082 3088 3102 3091
rect 3110 3091 3113 3098
rect 3750 3092 3753 3098
rect 3110 3088 3166 3091
rect 3258 3088 3350 3091
rect 3530 3088 3694 3091
rect 3706 3088 3718 3091
rect 582 3082 585 3088
rect 966 3082 969 3088
rect 1598 3082 1601 3088
rect 26 3078 46 3081
rect 50 3078 206 3081
rect 778 3078 782 3081
rect 802 3078 910 3081
rect 1058 3078 1134 3081
rect 1266 3078 1454 3081
rect 1474 3078 1574 3081
rect 1634 3078 1646 3081
rect 1658 3078 1662 3081
rect 1666 3078 1734 3081
rect 1738 3078 1934 3081
rect 2010 3078 2198 3081
rect 2202 3078 2270 3081
rect 2274 3078 2326 3081
rect 2330 3078 2494 3081
rect 2498 3078 2566 3081
rect 2578 3078 2654 3081
rect 2806 3078 2854 3081
rect 2858 3078 2974 3081
rect 3090 3078 3121 3081
rect 3186 3078 3198 3081
rect 3202 3078 3430 3081
rect 3538 3078 3614 3081
rect 3618 3078 3630 3081
rect 3658 3078 3678 3081
rect 3706 3078 3710 3081
rect 230 3072 233 3078
rect 566 3072 569 3078
rect 134 3068 214 3071
rect 450 3068 486 3071
rect 650 3068 734 3071
rect 738 3068 742 3071
rect 786 3068 854 3071
rect 858 3068 1078 3071
rect 1082 3068 1094 3071
rect 1098 3068 1110 3071
rect 1386 3068 1398 3071
rect 1410 3068 1478 3071
rect 1482 3068 1486 3071
rect 1538 3068 1670 3071
rect 1674 3068 1678 3071
rect 1690 3068 1710 3071
rect 1930 3068 1982 3071
rect 1986 3068 2014 3071
rect 2026 3068 2038 3071
rect 2042 3068 2214 3071
rect 2258 3068 2270 3071
rect 2402 3068 2438 3071
rect 2578 3068 2582 3071
rect 2670 3071 2673 3078
rect 2614 3068 2673 3071
rect 2806 3072 2809 3078
rect 3018 3068 3110 3071
rect 3118 3071 3121 3078
rect 3510 3072 3513 3078
rect 3118 3068 3206 3071
rect 3242 3068 3254 3071
rect 3298 3068 3310 3071
rect 3514 3068 3649 3071
rect 3666 3068 3742 3071
rect 134 3062 137 3068
rect 238 3062 241 3068
rect 2302 3062 2305 3068
rect 2614 3062 2617 3068
rect 226 3058 230 3061
rect 346 3058 670 3061
rect 746 3058 782 3061
rect 850 3058 950 3061
rect 1138 3058 1374 3061
rect 1378 3058 1422 3061
rect 1458 3058 1470 3061
rect 1506 3058 1526 3061
rect 1534 3058 1542 3061
rect 1546 3058 1550 3061
rect 1562 3058 1686 3061
rect 2002 3058 2006 3061
rect 2034 3058 2070 3061
rect 2074 3058 2134 3061
rect 2138 3058 2142 3061
rect 2162 3058 2166 3061
rect 2186 3058 2262 3061
rect 2274 3058 2278 3061
rect 2306 3058 2358 3061
rect 2430 3058 2438 3061
rect 2458 3058 2462 3061
rect 2570 3058 2590 3061
rect 2610 3058 2614 3061
rect 2674 3058 2694 3061
rect 2714 3058 2758 3061
rect 3066 3058 3070 3061
rect 3074 3058 3094 3061
rect 3130 3058 3142 3061
rect 3186 3058 3206 3061
rect 3210 3058 3238 3061
rect 3266 3058 3334 3061
rect 3474 3058 3478 3061
rect 3498 3058 3518 3061
rect 3626 3058 3630 3061
rect 3646 3061 3649 3068
rect 3646 3058 3742 3061
rect -26 3051 -22 3052
rect -26 3048 6 3051
rect 26 3048 246 3051
rect 458 3048 518 3051
rect 738 3048 806 3051
rect 818 3048 830 3051
rect 1010 3048 1086 3051
rect 1114 3048 1182 3051
rect 1242 3048 1326 3051
rect 1354 3048 1390 3051
rect 1394 3048 1398 3051
rect 1430 3051 1433 3058
rect 1430 3048 1494 3051
rect 1594 3048 1598 3051
rect 1642 3048 1670 3051
rect 1742 3051 1745 3058
rect 2422 3052 2425 3058
rect 2430 3052 2433 3058
rect 1678 3048 1745 3051
rect 1930 3048 1966 3051
rect 1970 3048 1982 3051
rect 1986 3048 2006 3051
rect 2042 3048 2062 3051
rect 2090 3048 2126 3051
rect 2130 3048 2230 3051
rect 2590 3051 2593 3058
rect 2462 3048 2481 3051
rect 2590 3048 2678 3051
rect 2882 3048 3118 3051
rect 3366 3051 3369 3058
rect 3234 3048 3430 3051
rect 3458 3048 3465 3051
rect 1678 3042 1681 3048
rect 1790 3042 1793 3048
rect 2462 3042 2465 3048
rect 2478 3042 2481 3048
rect 2694 3042 2697 3048
rect 234 3038 598 3041
rect 666 3038 670 3041
rect 770 3038 926 3041
rect 954 3038 1062 3041
rect 1082 3038 1134 3041
rect 1138 3038 1174 3041
rect 1394 3038 1425 3041
rect 1466 3038 1550 3041
rect 1626 3038 1630 3041
rect 1890 3038 2102 3041
rect 2122 3038 2134 3041
rect 2138 3038 2254 3041
rect 2274 3038 2366 3041
rect 2370 3038 2446 3041
rect 2570 3038 2598 3041
rect 2602 3038 2646 3041
rect 2650 3038 2654 3041
rect 3126 3041 3129 3048
rect 3462 3042 3465 3048
rect 3530 3048 3534 3051
rect 3570 3048 3582 3051
rect 3602 3048 3657 3051
rect 3666 3048 3694 3051
rect 3738 3048 3750 3051
rect 3058 3038 3238 3041
rect 3242 3038 3382 3041
rect 3402 3038 3406 3041
rect 3518 3041 3521 3048
rect 3590 3042 3593 3048
rect 3518 3038 3534 3041
rect 3654 3041 3657 3048
rect 3654 3038 3702 3041
rect 1422 3032 1425 3038
rect 362 3028 366 3031
rect 626 3028 902 3031
rect 1034 3028 1110 3031
rect 1122 3028 1174 3031
rect 1178 3028 1406 3031
rect 1450 3028 1606 3031
rect 1766 3031 1769 3038
rect 1766 3028 1926 3031
rect 1930 3028 2102 3031
rect 2114 3028 2126 3031
rect 2282 3028 2342 3031
rect 2346 3028 2382 3031
rect 2418 3028 2534 3031
rect 2542 3031 2545 3038
rect 2542 3028 2822 3031
rect 3290 3028 3518 3031
rect 506 3018 622 3021
rect 626 3018 1414 3021
rect 1418 3018 1430 3021
rect 1722 3018 1846 3021
rect 1930 3018 1998 3021
rect 2002 3018 2070 3021
rect 2082 3018 2270 3021
rect 2374 3018 2486 3021
rect 2530 3018 2878 3021
rect 3034 3018 3270 3021
rect 3274 3018 3326 3021
rect 3330 3018 3406 3021
rect 3418 3018 3454 3021
rect 3514 3018 3526 3021
rect 90 3008 118 3011
rect 586 3008 766 3011
rect 858 3008 862 3011
rect 866 3008 1126 3011
rect 2374 3011 2377 3018
rect 1522 3008 2377 3011
rect 2466 3008 2510 3011
rect 3026 3008 3062 3011
rect 3146 3008 3150 3011
rect 3298 3008 3310 3011
rect 3562 3008 3686 3011
rect 344 3003 346 3007
rect 350 3003 353 3007
rect 358 3003 360 3007
rect 1360 3003 1362 3007
rect 1366 3003 1369 3007
rect 1374 3003 1376 3007
rect 2384 3003 2386 3007
rect 2390 3003 2393 3007
rect 2398 3003 2400 3007
rect 3408 3003 3410 3007
rect 3414 3003 3417 3007
rect 3422 3003 3424 3007
rect 498 2998 694 3001
rect 698 2998 766 3001
rect 786 2998 894 3001
rect 922 2998 950 3001
rect 962 2998 1078 3001
rect 1394 2998 1574 3001
rect 1634 2998 1790 3001
rect 1794 2998 1878 3001
rect 2066 2998 2110 3001
rect 2130 2998 2334 3001
rect 2586 2998 2726 3001
rect 2730 2998 2750 3001
rect 3050 2998 3182 3001
rect 3186 2998 3401 3001
rect 3482 2998 3566 3001
rect 594 2988 598 2991
rect 782 2988 790 2991
rect 794 2988 918 2991
rect 922 2988 1262 2991
rect 1266 2988 1278 2991
rect 1282 2988 1542 2991
rect 1570 2988 1582 2991
rect 1666 2988 1782 2991
rect 1786 2988 1830 2991
rect 1962 2988 2238 2991
rect 2322 2988 3150 2991
rect 3274 2988 3334 2991
rect 3398 2991 3401 2998
rect 3398 2988 3446 2991
rect 3462 2988 3614 2991
rect 578 2978 638 2981
rect 658 2978 678 2981
rect 710 2981 713 2988
rect 3462 2982 3465 2988
rect 682 2978 713 2981
rect 762 2978 878 2981
rect 970 2978 1254 2981
rect 1262 2978 1270 2981
rect 1274 2978 1294 2981
rect 1330 2978 1446 2981
rect 1478 2978 1662 2981
rect 1666 2978 1670 2981
rect 2058 2978 2070 2981
rect 2106 2978 2201 2981
rect 2354 2978 2462 2981
rect 2466 2978 2502 2981
rect 2506 2978 2566 2981
rect 2618 2978 2622 2981
rect 2722 2978 3126 2981
rect 3138 2978 3337 2981
rect 3346 2978 3414 2981
rect 3522 2978 3590 2981
rect 1262 2972 1265 2978
rect 642 2968 694 2971
rect 714 2968 750 2971
rect 754 2968 814 2971
rect 818 2968 918 2971
rect 922 2968 1006 2971
rect 1010 2968 1046 2971
rect 1226 2968 1230 2971
rect 1318 2971 1321 2978
rect 1290 2968 1321 2971
rect 1478 2971 1481 2978
rect 1974 2972 1977 2978
rect 2030 2972 2033 2978
rect 2046 2972 2049 2978
rect 2054 2972 2057 2978
rect 1378 2968 1481 2971
rect 1490 2968 1550 2971
rect 1558 2968 1574 2971
rect 1610 2968 1622 2971
rect 1690 2968 1953 2971
rect 2010 2968 2014 2971
rect 2094 2971 2097 2978
rect 2198 2972 2201 2978
rect 2094 2968 2142 2971
rect 2146 2968 2190 2971
rect 2218 2968 2222 2971
rect 2266 2968 2326 2971
rect 2378 2968 2406 2971
rect 2458 2968 2478 2971
rect 2530 2968 2542 2971
rect 2554 2968 2982 2971
rect 3194 2968 3230 2971
rect 3258 2968 3270 2971
rect 3334 2971 3337 2978
rect 3334 2968 3350 2971
rect 3514 2968 3582 2971
rect 542 2961 545 2968
rect 522 2958 545 2961
rect 630 2961 633 2968
rect 1558 2962 1561 2968
rect 630 2958 649 2961
rect 754 2958 814 2961
rect 818 2958 870 2961
rect 914 2958 918 2961
rect 930 2958 942 2961
rect 946 2958 974 2961
rect 1210 2958 1230 2961
rect 1234 2958 1270 2961
rect 1290 2958 1310 2961
rect 1322 2958 1326 2961
rect 1458 2958 1470 2961
rect 1474 2958 1478 2961
rect 1618 2958 1678 2961
rect 1950 2961 1953 2968
rect 1950 2958 2270 2961
rect 2322 2958 2350 2961
rect 2430 2961 2433 2968
rect 3158 2962 3161 2968
rect 3318 2962 3321 2968
rect 2402 2958 2433 2961
rect 2458 2958 2462 2961
rect 2474 2958 2958 2961
rect 2978 2958 3126 2961
rect 3242 2958 3286 2961
rect 3322 2958 3390 2961
rect 3502 2961 3505 2968
rect 3498 2958 3534 2961
rect -26 2951 -22 2952
rect -26 2948 6 2951
rect 558 2951 561 2958
rect 558 2948 574 2951
rect 610 2948 614 2951
rect 646 2951 649 2958
rect 646 2948 830 2951
rect 842 2948 854 2951
rect 858 2948 942 2951
rect 946 2948 1689 2951
rect 1718 2951 1721 2958
rect 1698 2948 1721 2951
rect 1726 2952 1729 2958
rect 1942 2952 1945 2958
rect 3622 2952 3625 2958
rect 3654 2952 3657 2958
rect 1986 2948 2334 2951
rect 2374 2948 2382 2951
rect 2386 2948 2422 2951
rect 2450 2948 2462 2951
rect 2522 2948 2678 2951
rect 2930 2948 2966 2951
rect 3322 2948 3326 2951
rect 3330 2948 3334 2951
rect 3346 2948 3374 2951
rect 3386 2948 3390 2951
rect 3466 2948 3470 2951
rect 3546 2948 3606 2951
rect 3674 2948 3678 2951
rect 3762 2948 3766 2951
rect 550 2942 553 2948
rect 82 2938 94 2941
rect 98 2938 166 2941
rect 170 2938 238 2941
rect 322 2938 334 2941
rect 602 2938 766 2941
rect 818 2938 934 2941
rect 946 2938 974 2941
rect 1086 2938 1222 2941
rect 1242 2938 1246 2941
rect 1274 2938 1302 2941
rect 1442 2938 1446 2941
rect 1450 2938 1510 2941
rect 1522 2938 1526 2941
rect 1546 2938 1550 2941
rect 1594 2938 1598 2941
rect 1610 2938 1614 2941
rect 1686 2941 1689 2948
rect 1686 2938 1950 2941
rect 2002 2938 2006 2941
rect 2026 2938 2062 2941
rect 2130 2938 2134 2941
rect 2202 2938 2222 2941
rect 2250 2938 2382 2941
rect 2434 2938 2454 2941
rect 2498 2938 2502 2941
rect 2506 2938 2574 2941
rect 2714 2938 2742 2941
rect 2746 2938 2766 2941
rect 3230 2941 3233 2948
rect 3302 2942 3305 2948
rect 3230 2938 3270 2941
rect 3306 2938 3422 2941
rect 3514 2938 3622 2941
rect 3650 2938 3654 2941
rect 3658 2938 3662 2941
rect 3698 2938 3742 2941
rect 26 2928 238 2931
rect 414 2931 417 2938
rect 1086 2932 1089 2938
rect 1406 2932 1409 2938
rect 314 2928 417 2931
rect 538 2928 574 2931
rect 578 2928 670 2931
rect 690 2928 694 2931
rect 730 2928 750 2931
rect 762 2928 806 2931
rect 874 2928 902 2931
rect 978 2928 982 2931
rect 1194 2928 1230 2931
rect 1234 2928 1302 2931
rect 1422 2931 1425 2938
rect 2070 2932 2073 2938
rect 2662 2932 2665 2938
rect 1422 2928 1462 2931
rect 1466 2928 1622 2931
rect 1834 2928 1838 2931
rect 1850 2928 2006 2931
rect 2018 2928 2030 2931
rect 2138 2928 2142 2931
rect 2210 2928 2294 2931
rect 2306 2928 2342 2931
rect 2354 2928 2374 2931
rect 2386 2928 2470 2931
rect 2610 2928 2622 2931
rect 2666 2928 2774 2931
rect 2854 2931 2857 2938
rect 2778 2928 2857 2931
rect 3174 2932 3177 2938
rect 3758 2932 3761 2938
rect 3266 2928 3286 2931
rect 3290 2928 3454 2931
rect 3466 2928 3526 2931
rect 3554 2928 3574 2931
rect 3706 2928 3734 2931
rect 506 2918 574 2921
rect 630 2918 638 2921
rect 642 2918 646 2921
rect 890 2918 910 2921
rect 938 2918 1006 2921
rect 1010 2918 1054 2921
rect 1402 2918 1462 2921
rect 1514 2918 1534 2921
rect 1570 2918 1662 2921
rect 1670 2921 1673 2928
rect 1670 2918 1862 2921
rect 1882 2918 2158 2921
rect 2186 2918 2222 2921
rect 2226 2918 2262 2921
rect 2274 2918 2286 2921
rect 2314 2918 2486 2921
rect 2538 2918 2614 2921
rect 2762 2918 2870 2921
rect 2922 2918 2926 2921
rect 3154 2918 3310 2921
rect 3366 2918 3374 2921
rect 3378 2918 3382 2921
rect 3386 2918 3390 2921
rect 3570 2918 3646 2921
rect 3694 2921 3697 2928
rect 3674 2918 3750 2921
rect 34 2908 70 2911
rect 530 2908 630 2911
rect 954 2908 1110 2911
rect 1130 2908 1142 2911
rect 1330 2908 1518 2911
rect 1538 2908 1742 2911
rect 1746 2908 1870 2911
rect 1906 2908 2046 2911
rect 2066 2908 2078 2911
rect 2122 2908 2294 2911
rect 2322 2908 2342 2911
rect 2378 2908 2486 2911
rect 2610 2908 2662 2911
rect 2690 2908 2798 2911
rect 2802 2908 2878 2911
rect 3106 2908 3662 2911
rect 848 2903 850 2907
rect 854 2903 857 2907
rect 862 2903 864 2907
rect 1880 2903 1882 2907
rect 1886 2903 1889 2907
rect 1894 2903 1896 2907
rect 2904 2903 2906 2907
rect 2910 2903 2913 2907
rect 2918 2903 2920 2907
rect 338 2898 342 2901
rect 466 2898 750 2901
rect 786 2898 814 2901
rect 974 2898 1334 2901
rect 1354 2898 1366 2901
rect 1642 2898 1678 2901
rect 1698 2898 1702 2901
rect 1826 2898 1854 2901
rect 2042 2898 2046 2901
rect 2074 2898 2118 2901
rect 2162 2898 2542 2901
rect 2546 2898 2726 2901
rect 3218 2898 3278 2901
rect 3298 2898 3526 2901
rect 3530 2898 3558 2901
rect 570 2888 654 2891
rect 658 2888 665 2891
rect 698 2888 702 2891
rect 706 2888 718 2891
rect 974 2891 977 2898
rect 742 2888 977 2891
rect 986 2888 990 2891
rect 1002 2888 1182 2891
rect 1338 2888 2198 2891
rect 2230 2888 2366 2891
rect 2370 2888 2422 2891
rect 2458 2888 2766 2891
rect 2770 2888 2886 2891
rect 3170 2888 3198 2891
rect 3250 2888 3262 2891
rect 3362 2888 3470 2891
rect 3490 2888 3670 2891
rect 3754 2888 3766 2891
rect 30 2881 33 2888
rect -26 2878 33 2881
rect 94 2881 97 2888
rect 58 2878 118 2881
rect 742 2881 745 2888
rect 602 2878 750 2881
rect 778 2878 918 2881
rect 1314 2878 1478 2881
rect 1498 2878 1502 2881
rect 1514 2878 1750 2881
rect 1754 2878 1798 2881
rect 1874 2878 2022 2881
rect 2098 2878 2102 2881
rect 2230 2881 2233 2888
rect 2106 2878 2233 2881
rect 2242 2878 2286 2881
rect 2302 2878 2398 2881
rect 2402 2878 2414 2881
rect 2634 2878 2646 2881
rect 2810 2878 2814 2881
rect 2826 2878 2830 2881
rect 2902 2881 2905 2888
rect 3206 2882 3209 2888
rect 2902 2878 2926 2881
rect 3314 2878 3366 2881
rect 3546 2878 3574 2881
rect 3610 2878 3654 2881
rect 3658 2878 3662 2881
rect 3706 2878 3734 2881
rect 3738 2878 3758 2881
rect -26 2872 -23 2878
rect 230 2872 233 2878
rect 1094 2872 1097 2878
rect 2302 2872 2305 2878
rect 2694 2872 2697 2878
rect -26 2868 -22 2872
rect 18 2868 206 2871
rect 458 2868 478 2871
rect 682 2868 750 2871
rect 754 2868 777 2871
rect 818 2868 822 2871
rect 858 2868 862 2871
rect 1186 2868 1206 2871
rect 1274 2868 1286 2871
rect 1290 2868 1294 2871
rect 1306 2868 1358 2871
rect 1370 2868 1430 2871
rect 1474 2868 1478 2871
rect 1698 2868 1702 2871
rect 1730 2868 1782 2871
rect 1786 2868 1982 2871
rect 1986 2868 2014 2871
rect 2026 2868 2102 2871
rect 2138 2868 2153 2871
rect 2162 2868 2198 2871
rect 2202 2868 2230 2871
rect 2338 2868 2342 2871
rect 2354 2868 2422 2871
rect 2474 2868 2614 2871
rect 2618 2868 2622 2871
rect 2754 2868 2758 2871
rect 2814 2871 2817 2878
rect 2814 2868 3054 2871
rect 3150 2871 3153 2878
rect 3114 2868 3153 2871
rect 3198 2868 3254 2871
rect 3282 2868 3334 2871
rect 3518 2871 3521 2878
rect 3426 2868 3521 2871
rect 3570 2868 3574 2871
rect 3626 2868 3630 2871
rect 774 2862 777 2868
rect 2150 2862 2153 2868
rect 3198 2862 3201 2868
rect 34 2858 38 2861
rect 58 2858 62 2861
rect 66 2858 118 2861
rect 122 2858 214 2861
rect 378 2858 422 2861
rect 426 2858 454 2861
rect 514 2858 686 2861
rect 762 2858 766 2861
rect 794 2858 822 2861
rect 842 2858 862 2861
rect 866 2858 886 2861
rect 914 2858 1070 2861
rect 1082 2858 1166 2861
rect 1186 2858 1422 2861
rect 1450 2858 1558 2861
rect 1626 2858 1766 2861
rect 1906 2858 1985 2861
rect 2018 2858 2038 2861
rect 2066 2858 2070 2861
rect 2082 2858 2086 2861
rect 2098 2858 2126 2861
rect 2138 2858 2142 2861
rect 2170 2858 2174 2861
rect 2210 2858 2214 2861
rect 2226 2858 2246 2861
rect 2386 2858 2390 2861
rect 2394 2858 2438 2861
rect 2578 2858 2582 2861
rect 2590 2858 2630 2861
rect 2634 2858 2638 2861
rect 2786 2858 2814 2861
rect 2994 2858 3086 2861
rect 3122 2858 3153 2861
rect 3266 2858 3382 2861
rect 3442 2858 3614 2861
rect 3690 2858 3726 2861
rect 1982 2852 1985 2858
rect 2278 2852 2281 2858
rect 2302 2852 2305 2858
rect 2590 2852 2593 2858
rect 2662 2852 2665 2858
rect 2710 2852 2713 2858
rect 3150 2852 3153 2858
rect -26 2851 -22 2852
rect -26 2848 6 2851
rect 50 2848 65 2851
rect 62 2842 65 2848
rect 130 2848 134 2851
rect 250 2848 254 2851
rect 602 2848 614 2851
rect 618 2848 854 2851
rect 858 2848 950 2851
rect 1202 2848 1334 2851
rect 1354 2848 1366 2851
rect 1474 2848 1606 2851
rect 1642 2848 1854 2851
rect 2082 2848 2254 2851
rect 2314 2848 2318 2851
rect 2362 2848 2518 2851
rect 2546 2848 2550 2851
rect 2602 2848 2622 2851
rect 2650 2848 2654 2851
rect 2690 2848 2694 2851
rect 2730 2848 3014 2851
rect 3042 2848 3046 2851
rect 3074 2848 3102 2851
rect 3294 2848 3302 2851
rect 3306 2848 3334 2851
rect 3346 2848 3350 2851
rect 3394 2848 3454 2851
rect 110 2842 113 2848
rect 570 2838 678 2841
rect 714 2838 718 2841
rect 730 2838 785 2841
rect 842 2838 870 2841
rect 874 2838 1006 2841
rect 1082 2838 1086 2841
rect 1090 2838 1270 2841
rect 1338 2838 1398 2841
rect 1474 2838 1486 2841
rect 1762 2838 1942 2841
rect 1978 2838 2198 2841
rect 2202 2838 2334 2841
rect 2346 2838 2502 2841
rect 2506 2838 2598 2841
rect 2722 2838 2990 2841
rect 3034 2838 3062 2841
rect 3066 2838 3094 2841
rect 3590 2841 3593 2848
rect 3098 2838 3593 2841
rect 782 2832 785 2838
rect 1046 2832 1049 2838
rect 162 2828 230 2831
rect 322 2828 742 2831
rect 1346 2828 1390 2831
rect 1410 2828 1454 2831
rect 1530 2828 1574 2831
rect 1746 2828 2462 2831
rect 2466 2828 2694 2831
rect 3042 2828 3070 2831
rect 3234 2828 3302 2831
rect 3306 2828 3318 2831
rect 3322 2828 3358 2831
rect 3366 2828 3398 2831
rect 3402 2828 3406 2831
rect 3418 2828 3550 2831
rect 3554 2828 3630 2831
rect 3366 2822 3369 2828
rect 74 2818 166 2821
rect 802 2818 878 2821
rect 898 2818 966 2821
rect 970 2818 1070 2821
rect 1298 2818 1798 2821
rect 1946 2818 1998 2821
rect 2002 2818 2150 2821
rect 2154 2818 2166 2821
rect 2226 2818 2446 2821
rect 2522 2818 2646 2821
rect 3498 2818 3542 2821
rect 90 2808 294 2811
rect 418 2808 550 2811
rect 690 2808 854 2811
rect 898 2808 1014 2811
rect 1026 2808 1046 2811
rect 1322 2808 1350 2811
rect 1386 2808 1518 2811
rect 1522 2808 1742 2811
rect 1762 2808 1766 2811
rect 1994 2808 2078 2811
rect 2098 2808 2102 2811
rect 2146 2808 2222 2811
rect 2258 2808 2342 2811
rect 2442 2808 2462 2811
rect 2538 2808 2862 2811
rect 2922 2808 2934 2811
rect 3746 2808 3774 2811
rect 344 2803 346 2807
rect 350 2803 353 2807
rect 358 2803 360 2807
rect 1360 2803 1362 2807
rect 1366 2803 1369 2807
rect 1374 2803 1376 2807
rect 2384 2803 2386 2807
rect 2390 2803 2393 2807
rect 2398 2803 2400 2807
rect 3408 2803 3410 2807
rect 3414 2803 3417 2807
rect 3422 2803 3424 2807
rect 58 2798 94 2801
rect 146 2798 214 2801
rect 658 2798 662 2801
rect 666 2798 806 2801
rect 810 2798 1302 2801
rect 1458 2798 1678 2801
rect 1682 2798 1758 2801
rect 1770 2798 1846 2801
rect 1858 2798 2374 2801
rect 2682 2798 2686 2801
rect 3130 2798 3158 2801
rect 3434 2798 3494 2801
rect 666 2788 777 2791
rect 646 2781 649 2788
rect 774 2782 777 2788
rect 890 2788 918 2791
rect 1130 2788 1134 2791
rect 1154 2788 1486 2791
rect 1738 2788 1790 2791
rect 1826 2788 1838 2791
rect 1842 2788 2006 2791
rect 2010 2788 2118 2791
rect 2122 2788 2254 2791
rect 2258 2788 2286 2791
rect 2290 2788 2390 2791
rect 2394 2788 2478 2791
rect 2634 2788 2734 2791
rect 2738 2788 2774 2791
rect 2914 2788 2918 2791
rect 3002 2788 3238 2791
rect 3442 2788 3446 2791
rect 806 2782 809 2788
rect 466 2778 649 2781
rect 714 2778 734 2781
rect 814 2778 929 2781
rect 1114 2778 1526 2781
rect 2170 2778 2238 2781
rect 2306 2778 3238 2781
rect 3438 2778 3566 2781
rect 3570 2778 3598 2781
rect 546 2768 550 2771
rect 554 2768 614 2771
rect 618 2768 718 2771
rect 762 2768 766 2771
rect 786 2768 790 2771
rect 798 2771 801 2778
rect 794 2768 801 2771
rect 814 2771 817 2778
rect 926 2772 929 2778
rect 810 2768 817 2771
rect 942 2768 1334 2771
rect 1418 2768 1422 2771
rect 1426 2768 1470 2771
rect 1710 2771 1713 2778
rect 3438 2772 3441 2778
rect 1710 2768 1726 2771
rect 1938 2768 1982 2771
rect 1986 2768 1993 2771
rect 2266 2768 2278 2771
rect 2290 2768 2318 2771
rect 2354 2768 2558 2771
rect 2562 2768 2630 2771
rect 2722 2768 2726 2771
rect 2794 2768 2798 2771
rect 3082 2768 3086 2771
rect 3202 2768 3294 2771
rect 3354 2768 3382 2771
rect 3538 2768 3558 2771
rect 3726 2771 3729 2778
rect 3722 2768 3729 2771
rect 3746 2768 3750 2771
rect 618 2758 622 2761
rect 714 2758 774 2761
rect 778 2758 790 2761
rect 838 2761 841 2768
rect 942 2762 945 2768
rect 798 2758 841 2761
rect 906 2758 926 2761
rect 1010 2758 1014 2761
rect 1034 2758 1054 2761
rect 1066 2758 1110 2761
rect 1250 2758 1366 2761
rect 1402 2758 1478 2761
rect 1618 2758 1622 2761
rect 1782 2761 1785 2768
rect 3518 2762 3521 2768
rect 1738 2758 1785 2761
rect 1858 2758 1902 2761
rect 1994 2758 2014 2761
rect 2026 2758 2118 2761
rect 2274 2758 2286 2761
rect 2314 2758 2334 2761
rect 2350 2758 2366 2761
rect 2458 2758 2478 2761
rect 2610 2758 2614 2761
rect 2666 2758 2742 2761
rect 2746 2758 2862 2761
rect 3178 2758 3270 2761
rect 3274 2758 3358 2761
rect 3458 2758 3502 2761
rect 3546 2758 3654 2761
rect 3666 2758 3686 2761
rect -26 2751 -22 2752
rect -26 2748 6 2751
rect 342 2751 345 2758
rect 338 2748 345 2751
rect 618 2748 710 2751
rect 798 2751 801 2758
rect 786 2748 801 2751
rect 826 2748 894 2751
rect 922 2748 1342 2751
rect 1402 2748 1438 2751
rect 1442 2748 1462 2751
rect 1466 2748 1678 2751
rect 1682 2748 1694 2751
rect 1702 2751 1705 2758
rect 1726 2751 1729 2758
rect 1702 2748 1729 2751
rect 1746 2748 1750 2751
rect 1818 2748 1849 2751
rect 1874 2748 1894 2751
rect 1986 2748 1990 2751
rect 2018 2748 2054 2751
rect 2178 2748 2270 2751
rect 2350 2751 2353 2758
rect 2346 2748 2353 2751
rect 2362 2748 2366 2751
rect 2378 2748 2542 2751
rect 2674 2748 2710 2751
rect 2714 2748 2782 2751
rect 2846 2748 2854 2751
rect 2858 2748 2878 2751
rect 2922 2748 3022 2751
rect 3082 2748 3086 2751
rect 3090 2748 3102 2751
rect 3274 2748 3278 2751
rect 3378 2748 3550 2751
rect 3554 2748 3590 2751
rect 3594 2748 3622 2751
rect 3658 2748 3673 2751
rect 3714 2748 3758 2751
rect 134 2742 137 2748
rect 310 2741 313 2748
rect 1846 2742 1849 2748
rect 310 2738 374 2741
rect 482 2738 526 2741
rect 570 2738 622 2741
rect 642 2738 726 2741
rect 746 2738 822 2741
rect 842 2738 846 2741
rect 890 2738 902 2741
rect 906 2738 910 2741
rect 914 2738 942 2741
rect 954 2738 958 2741
rect 978 2738 1030 2741
rect 1034 2738 1062 2741
rect 1066 2738 1094 2741
rect 1346 2738 1406 2741
rect 1458 2738 1486 2741
rect 1490 2738 1550 2741
rect 1554 2738 1686 2741
rect 1690 2738 1702 2741
rect 1746 2738 1809 2741
rect 1890 2738 1942 2741
rect 1946 2738 2022 2741
rect 2034 2738 2049 2741
rect 2098 2738 2246 2741
rect 2294 2741 2297 2748
rect 3670 2742 3673 2748
rect 2250 2738 2297 2741
rect 2378 2738 2422 2741
rect 2450 2738 2470 2741
rect 2638 2738 2646 2741
rect 2650 2738 2662 2741
rect 2690 2738 2766 2741
rect 2794 2738 2798 2741
rect 2826 2738 2846 2741
rect 3266 2738 3422 2741
rect 3474 2738 3502 2741
rect 3506 2738 3614 2741
rect 3618 2738 3622 2741
rect 3626 2738 3646 2741
rect 478 2731 481 2738
rect 298 2728 481 2731
rect 638 2732 641 2738
rect 1214 2732 1217 2738
rect 1230 2732 1233 2738
rect 1438 2732 1441 2738
rect 1806 2732 1809 2738
rect 2046 2732 2049 2738
rect 666 2728 670 2731
rect 714 2728 830 2731
rect 882 2728 934 2731
rect 954 2728 990 2731
rect 1018 2728 1022 2731
rect 1514 2728 1646 2731
rect 1674 2728 1694 2731
rect 1818 2728 1910 2731
rect 1954 2728 1958 2731
rect 2210 2728 2286 2731
rect 2402 2728 2454 2731
rect 2458 2728 2478 2731
rect 2562 2728 2734 2731
rect 2778 2728 2830 2731
rect 3006 2731 3009 2738
rect 2930 2728 3009 2731
rect 3362 2728 3414 2731
rect 3470 2731 3473 2738
rect 3418 2728 3473 2731
rect 3530 2728 3534 2731
rect 3578 2728 3742 2731
rect 3746 2728 3774 2731
rect 426 2718 902 2721
rect 906 2718 998 2721
rect 1046 2721 1049 2728
rect 2038 2722 2041 2728
rect 1046 2718 1062 2721
rect 1122 2718 1294 2721
rect 1414 2718 1526 2721
rect 1530 2718 1590 2721
rect 1690 2718 1734 2721
rect 1858 2718 1910 2721
rect 1978 2718 1982 2721
rect 2074 2718 2406 2721
rect 2442 2718 2598 2721
rect 2642 2718 2654 2721
rect 2818 2718 3174 2721
rect 3282 2718 3326 2721
rect 3398 2718 3406 2721
rect 3410 2718 3518 2721
rect 3530 2718 3614 2721
rect 3618 2718 3638 2721
rect 3650 2718 3678 2721
rect 3722 2718 3734 2721
rect 3738 2718 3750 2721
rect 82 2708 214 2711
rect 218 2708 318 2711
rect 402 2708 478 2711
rect 522 2708 670 2711
rect 834 2708 838 2711
rect 898 2708 958 2711
rect 970 2708 1038 2711
rect 1414 2711 1417 2718
rect 1050 2708 1417 2711
rect 1426 2708 1702 2711
rect 1722 2708 1726 2711
rect 1786 2708 1862 2711
rect 1906 2708 2022 2711
rect 2026 2708 2110 2711
rect 2138 2708 2142 2711
rect 2210 2708 2214 2711
rect 2250 2708 2366 2711
rect 2370 2708 2398 2711
rect 2418 2708 2494 2711
rect 2962 2708 3262 2711
rect 3290 2708 3294 2711
rect 3338 2708 3374 2711
rect 3402 2708 3542 2711
rect 3546 2708 3710 2711
rect 848 2703 850 2707
rect 854 2703 857 2707
rect 862 2703 864 2707
rect 1880 2703 1882 2707
rect 1886 2703 1889 2707
rect 1894 2703 1896 2707
rect 2702 2702 2705 2708
rect 2774 2702 2777 2708
rect 2904 2703 2906 2707
rect 2910 2703 2913 2707
rect 2918 2703 2920 2707
rect 634 2698 710 2701
rect 930 2698 1078 2701
rect 1082 2698 1350 2701
rect 1354 2698 1494 2701
rect 1634 2698 1790 2701
rect 1794 2698 1862 2701
rect 1866 2698 1870 2701
rect 1922 2698 2110 2701
rect 2450 2698 2462 2701
rect 2466 2698 2630 2701
rect 2634 2698 2646 2701
rect 2682 2698 2694 2701
rect 2858 2698 2862 2701
rect 3058 2698 3142 2701
rect 3170 2698 3350 2701
rect 3490 2698 3526 2701
rect 3546 2698 3558 2701
rect 3586 2698 3670 2701
rect 878 2692 881 2698
rect 894 2692 897 2698
rect 466 2688 582 2691
rect 586 2688 598 2691
rect 610 2688 774 2691
rect 850 2688 870 2691
rect 922 2688 950 2691
rect 978 2688 998 2691
rect 1034 2688 1126 2691
rect 1146 2688 1150 2691
rect 1154 2688 1166 2691
rect 1482 2688 1494 2691
rect 1498 2688 1534 2691
rect 1638 2688 1646 2691
rect 1650 2688 1662 2691
rect 1674 2688 1726 2691
rect 1762 2688 2078 2691
rect 2250 2688 2422 2691
rect 2426 2688 2446 2691
rect 2642 2688 2934 2691
rect 3266 2688 3486 2691
rect 3546 2688 3566 2691
rect 3626 2688 3630 2691
rect 366 2681 369 2688
rect 366 2678 422 2681
rect 570 2678 590 2681
rect 634 2678 758 2681
rect 770 2678 782 2681
rect 802 2678 806 2681
rect 866 2678 926 2681
rect 986 2678 990 2681
rect 1082 2678 1086 2681
rect 1130 2678 1310 2681
rect 1566 2681 1569 2688
rect 3046 2682 3049 2688
rect 1394 2678 1569 2681
rect 1578 2678 1678 2681
rect 1698 2678 1942 2681
rect 1994 2678 2158 2681
rect 2226 2678 2238 2681
rect 2274 2678 2350 2681
rect 2418 2678 2646 2681
rect 2654 2678 2718 2681
rect 2722 2678 3046 2681
rect 3122 2678 3166 2681
rect 3186 2678 3190 2681
rect 3194 2678 3294 2681
rect 3590 2681 3593 2688
rect 3298 2678 3593 2681
rect 3658 2678 3694 2681
rect 10 2668 70 2671
rect 214 2671 217 2678
rect 214 2668 406 2671
rect 430 2671 433 2678
rect 1998 2672 2001 2678
rect 2254 2672 2257 2678
rect 2366 2672 2369 2678
rect 430 2668 630 2671
rect 642 2668 646 2671
rect 730 2668 734 2671
rect 754 2668 958 2671
rect 962 2668 1014 2671
rect 1082 2668 1086 2671
rect 1106 2668 1222 2671
rect 1226 2668 1406 2671
rect 1450 2668 1558 2671
rect 1586 2668 1590 2671
rect 1618 2668 1654 2671
rect 1690 2668 1718 2671
rect 1722 2668 1742 2671
rect 1802 2668 1838 2671
rect 1842 2668 1878 2671
rect 1930 2668 1958 2671
rect 2122 2668 2134 2671
rect 2162 2668 2166 2671
rect 2194 2668 2214 2671
rect 2234 2668 2246 2671
rect 2262 2668 2342 2671
rect 2382 2668 2446 2671
rect 2654 2671 2657 2678
rect 2546 2668 2657 2671
rect 2682 2668 2686 2671
rect 2698 2668 2702 2671
rect 2738 2668 2798 2671
rect 2818 2668 2838 2671
rect 2850 2668 2854 2671
rect 2858 2668 2862 2671
rect 2898 2668 2902 2671
rect 2930 2668 2942 2671
rect 3162 2668 3198 2671
rect 3202 2668 3214 2671
rect 3218 2668 3222 2671
rect 3226 2668 3278 2671
rect 3282 2668 3286 2671
rect 3330 2668 3510 2671
rect 3530 2668 3606 2671
rect 3610 2668 3630 2671
rect 1038 2662 1041 2668
rect 322 2658 334 2661
rect 338 2658 342 2661
rect 362 2658 382 2661
rect 402 2658 454 2661
rect 458 2658 462 2661
rect 514 2658 542 2661
rect 546 2658 574 2661
rect 706 2658 918 2661
rect 946 2658 950 2661
rect 978 2658 1022 2661
rect 1242 2658 1246 2661
rect 1298 2658 1334 2661
rect 1562 2658 1638 2661
rect 1642 2658 1758 2661
rect 1762 2658 1766 2661
rect 1834 2658 2086 2661
rect 2146 2658 2150 2661
rect 2262 2661 2265 2668
rect 2250 2658 2265 2661
rect 2382 2661 2385 2668
rect 2322 2658 2385 2661
rect 2418 2658 2598 2661
rect 2654 2658 2726 2661
rect 2730 2658 2878 2661
rect 2886 2661 2889 2668
rect 2886 2658 3030 2661
rect 3186 2658 3190 2661
rect 3218 2658 3654 2661
rect 3714 2658 3726 2661
rect 502 2652 505 2658
rect -26 2651 -22 2652
rect -26 2648 366 2651
rect 378 2648 382 2651
rect 418 2648 489 2651
rect 586 2648 590 2651
rect 702 2651 705 2658
rect 626 2648 705 2651
rect 722 2648 742 2651
rect 882 2648 902 2651
rect 914 2648 1198 2651
rect 1226 2648 1302 2651
rect 1510 2651 1513 2658
rect 1806 2652 1809 2658
rect 1822 2652 1825 2658
rect 2654 2652 2657 2658
rect 1510 2648 1702 2651
rect 1706 2648 1726 2651
rect 1738 2648 1782 2651
rect 1842 2648 2110 2651
rect 2266 2648 2278 2651
rect 2386 2648 2406 2651
rect 2418 2648 2422 2651
rect 2450 2648 2654 2651
rect 2666 2648 2718 2651
rect 2722 2648 2846 2651
rect 2866 2648 2966 2651
rect 2970 2648 3078 2651
rect 3098 2648 3198 2651
rect 3234 2648 3334 2651
rect 3346 2648 3382 2651
rect 3426 2648 3470 2651
rect 3498 2648 3510 2651
rect 3538 2648 3550 2651
rect 3570 2648 3622 2651
rect 3714 2648 3774 2651
rect 486 2642 489 2648
rect 3654 2642 3657 2648
rect 474 2638 478 2641
rect 506 2638 558 2641
rect 578 2638 686 2641
rect 698 2638 718 2641
rect 738 2638 758 2641
rect 778 2638 1182 2641
rect 1298 2638 2214 2641
rect 2298 2638 2502 2641
rect 2506 2638 2654 2641
rect 2754 2638 2758 2641
rect 2774 2638 2798 2641
rect 2826 2638 2830 2641
rect 2842 2638 2854 2641
rect 2906 2638 3062 2641
rect 3066 2638 3118 2641
rect 3250 2638 3566 2641
rect 3578 2638 3590 2641
rect 446 2631 449 2638
rect 446 2628 734 2631
rect 794 2628 830 2631
rect 834 2628 846 2631
rect 898 2628 918 2631
rect 986 2628 990 2631
rect 1018 2628 1086 2631
rect 1106 2628 1153 2631
rect 1258 2628 1598 2631
rect 1666 2628 1734 2631
rect 1754 2628 1814 2631
rect 1818 2628 1934 2631
rect 1946 2628 1958 2631
rect 2018 2628 2294 2631
rect 2298 2628 2305 2631
rect 2314 2628 2406 2631
rect 2670 2631 2673 2638
rect 2562 2628 2673 2631
rect 2742 2632 2745 2638
rect 2774 2632 2777 2638
rect 2810 2628 2862 2631
rect 3194 2628 3406 2631
rect 3506 2628 3726 2631
rect 1006 2622 1009 2628
rect 650 2618 766 2621
rect 770 2618 806 2621
rect 810 2618 982 2621
rect 1010 2618 1142 2621
rect 1150 2621 1153 2628
rect 1150 2618 1286 2621
rect 1554 2618 1582 2621
rect 1610 2618 1926 2621
rect 1930 2618 2278 2621
rect 2282 2618 2721 2621
rect 2794 2618 3094 2621
rect 3106 2618 3230 2621
rect 3266 2618 3454 2621
rect 370 2608 846 2611
rect 906 2608 918 2611
rect 1066 2608 1294 2611
rect 1586 2608 1662 2611
rect 1730 2608 1862 2611
rect 1898 2608 1918 2611
rect 1922 2608 1942 2611
rect 2098 2608 2206 2611
rect 2282 2608 2374 2611
rect 2410 2608 2542 2611
rect 2718 2611 2721 2618
rect 2546 2608 2681 2611
rect 2718 2608 2998 2611
rect 3258 2608 3374 2611
rect 3506 2608 3598 2611
rect 344 2603 346 2607
rect 350 2603 353 2607
rect 358 2603 360 2607
rect 1046 2602 1049 2608
rect 1360 2603 1362 2607
rect 1366 2603 1369 2607
rect 1374 2603 1376 2607
rect 2384 2603 2386 2607
rect 2390 2603 2393 2607
rect 2398 2603 2400 2607
rect 602 2598 862 2601
rect 874 2598 894 2601
rect 898 2598 974 2601
rect 1082 2598 1246 2601
rect 1482 2598 1542 2601
rect 1590 2598 1614 2601
rect 1618 2598 2158 2601
rect 2162 2598 2377 2601
rect 2410 2598 2534 2601
rect 2554 2598 2670 2601
rect 2678 2601 2681 2608
rect 3408 2603 3410 2607
rect 3414 2603 3417 2607
rect 3422 2603 3424 2607
rect 2678 2598 2990 2601
rect 2994 2598 3398 2601
rect 3498 2598 3670 2601
rect 394 2588 782 2591
rect 802 2588 830 2591
rect 842 2588 926 2591
rect 1590 2591 1593 2598
rect 978 2588 1593 2591
rect 1602 2588 1798 2591
rect 1802 2588 2294 2591
rect 2306 2588 2318 2591
rect 2374 2591 2377 2598
rect 2374 2588 2710 2591
rect 2714 2588 2838 2591
rect 2858 2588 2942 2591
rect 3210 2588 3526 2591
rect 122 2578 142 2581
rect 658 2578 670 2581
rect 934 2581 937 2588
rect 674 2578 958 2581
rect 962 2578 1118 2581
rect 1154 2578 1502 2581
rect 1754 2578 1950 2581
rect 1954 2578 2246 2581
rect 2266 2578 2390 2581
rect 2466 2578 2585 2581
rect 2602 2578 2702 2581
rect 2818 2578 2830 2581
rect 2834 2578 2838 2581
rect 2898 2578 2958 2581
rect 3050 2578 3086 2581
rect 3090 2578 3110 2581
rect 3114 2578 3214 2581
rect 3218 2578 3254 2581
rect 3418 2578 3526 2581
rect 3594 2578 3646 2581
rect 3650 2578 3702 2581
rect 1518 2572 1521 2578
rect 2582 2572 2585 2578
rect 2782 2572 2785 2578
rect 714 2568 758 2571
rect 762 2568 766 2571
rect 770 2568 822 2571
rect 890 2568 894 2571
rect 954 2568 974 2571
rect 1058 2568 1150 2571
rect 1178 2568 1206 2571
rect 1346 2568 1390 2571
rect 1790 2568 1806 2571
rect 2122 2568 2134 2571
rect 2138 2568 2422 2571
rect 2718 2568 2758 2571
rect 2790 2571 2793 2578
rect 2790 2568 2830 2571
rect 2890 2568 3070 2571
rect 3074 2568 3174 2571
rect 3182 2568 3318 2571
rect 3330 2568 3334 2571
rect 3442 2568 3478 2571
rect 3602 2568 3614 2571
rect 646 2562 649 2568
rect 654 2562 657 2568
rect -26 2561 -22 2562
rect -26 2558 6 2561
rect 674 2558 694 2561
rect 722 2558 726 2561
rect 762 2558 798 2561
rect 898 2558 902 2561
rect 1006 2561 1009 2568
rect 1790 2562 1793 2568
rect 914 2558 1009 2561
rect 1082 2558 1270 2561
rect 1274 2558 1278 2561
rect 1522 2558 1758 2561
rect 1770 2558 1774 2561
rect 1834 2558 1838 2561
rect 1898 2558 1910 2561
rect 2122 2558 2145 2561
rect 2154 2558 2374 2561
rect 2386 2558 2454 2561
rect 2466 2558 2494 2561
rect 2506 2558 2510 2561
rect 2550 2561 2553 2568
rect 2538 2558 2553 2561
rect 2718 2562 2721 2568
rect 2862 2562 2865 2568
rect 3182 2562 3185 2568
rect 2794 2558 2798 2561
rect 2842 2558 2846 2561
rect 2874 2558 2974 2561
rect 3042 2558 3174 2561
rect 3210 2558 3222 2561
rect 3234 2558 3238 2561
rect 3266 2558 3342 2561
rect 3346 2558 3350 2561
rect 3354 2558 3470 2561
rect 3474 2558 3550 2561
rect 3590 2561 3593 2568
rect 3554 2558 3606 2561
rect 3614 2558 3686 2561
rect 3694 2561 3697 2568
rect 3758 2561 3761 2568
rect 3694 2558 3761 2561
rect 1382 2552 1385 2558
rect 2142 2552 2145 2558
rect 3614 2552 3617 2558
rect 138 2548 158 2551
rect 370 2548 446 2551
rect 682 2548 694 2551
rect 698 2548 742 2551
rect 746 2548 798 2551
rect 802 2548 806 2551
rect 834 2548 878 2551
rect 954 2548 982 2551
rect 986 2548 1094 2551
rect 1126 2548 1230 2551
rect 1386 2548 1574 2551
rect 1634 2548 1774 2551
rect 1798 2548 1806 2551
rect 1818 2548 1822 2551
rect 1914 2548 1934 2551
rect 1962 2548 1974 2551
rect 2170 2548 2326 2551
rect 2330 2548 2430 2551
rect 2434 2548 2502 2551
rect 2506 2548 2582 2551
rect 2602 2548 2614 2551
rect 2658 2548 2662 2551
rect 2690 2548 2710 2551
rect 2738 2548 2982 2551
rect 3002 2548 3030 2551
rect 3066 2548 3166 2551
rect 3178 2548 3326 2551
rect 3402 2548 3494 2551
rect 3506 2548 3510 2551
rect 3522 2548 3542 2551
rect 3642 2548 3662 2551
rect 3770 2548 3822 2551
rect -26 2538 -22 2542
rect 186 2538 254 2541
rect 502 2541 505 2548
rect 1126 2542 1129 2548
rect 2118 2542 2121 2548
rect 502 2538 574 2541
rect 634 2538 734 2541
rect 738 2538 758 2541
rect 850 2538 878 2541
rect 890 2538 894 2541
rect 922 2538 974 2541
rect 1098 2538 1102 2541
rect 1138 2538 1142 2541
rect 1178 2538 1182 2541
rect 1202 2538 1246 2541
rect 1266 2538 1478 2541
rect 1506 2538 1510 2541
rect 1554 2538 1694 2541
rect 1738 2538 1766 2541
rect 1786 2538 1798 2541
rect 1850 2538 1902 2541
rect 1978 2538 2102 2541
rect 2122 2538 2166 2541
rect 2186 2538 2342 2541
rect 2346 2538 2462 2541
rect 2474 2538 2510 2541
rect 2514 2538 2742 2541
rect 2754 2538 2774 2541
rect 2810 2538 2886 2541
rect 2898 2538 2902 2541
rect 3098 2538 3118 2541
rect 3130 2538 3222 2541
rect 3226 2538 3254 2541
rect 3370 2538 3446 2541
rect 3518 2541 3521 2548
rect 3450 2538 3521 2541
rect 3614 2542 3617 2548
rect 3650 2538 3678 2541
rect 3738 2538 3742 2541
rect 294 2531 297 2538
rect 1126 2532 1129 2538
rect 82 2528 297 2531
rect 386 2528 414 2531
rect 418 2528 606 2531
rect 786 2528 918 2531
rect 946 2528 1062 2531
rect 1066 2528 1102 2531
rect 1218 2528 1222 2531
rect 1234 2528 1270 2531
rect 1290 2528 1542 2531
rect 1626 2528 1649 2531
rect 1666 2528 1849 2531
rect 2098 2528 2142 2531
rect 2146 2528 2150 2531
rect 2266 2528 2302 2531
rect 2322 2528 2334 2531
rect 2410 2528 2574 2531
rect 2602 2528 2638 2531
rect 2802 2528 2822 2531
rect 2858 2528 2862 2531
rect 2890 2528 2942 2531
rect 3018 2528 3070 2531
rect 3074 2528 3102 2531
rect 3106 2528 3150 2531
rect 3154 2528 3214 2531
rect 3218 2528 3278 2531
rect 3386 2528 3398 2531
rect 3410 2528 3454 2531
rect 1646 2522 1649 2528
rect 1846 2522 1849 2528
rect 2246 2522 2249 2528
rect 3494 2522 3497 2528
rect 122 2518 174 2521
rect 218 2518 222 2521
rect 562 2518 710 2521
rect 714 2518 782 2521
rect 810 2518 822 2521
rect 826 2518 1078 2521
rect 1130 2518 1158 2521
rect 1162 2518 1198 2521
rect 1210 2518 1342 2521
rect 1346 2518 1550 2521
rect 1786 2518 1822 2521
rect 1866 2518 1982 2521
rect 2082 2518 2182 2521
rect 2338 2518 2390 2521
rect 2426 2518 2438 2521
rect 2514 2518 2542 2521
rect 2610 2518 2630 2521
rect 2882 2518 3094 2521
rect 3122 2518 3134 2521
rect 3226 2518 3262 2521
rect 3578 2518 3646 2521
rect 130 2508 134 2511
rect 466 2508 478 2511
rect 482 2508 622 2511
rect 690 2508 750 2511
rect 754 2508 782 2511
rect 786 2508 814 2511
rect 874 2508 958 2511
rect 986 2508 1062 2511
rect 1098 2508 1190 2511
rect 1234 2508 1238 2511
rect 1290 2508 1542 2511
rect 1570 2508 1662 2511
rect 1666 2508 1782 2511
rect 1794 2508 1838 2511
rect 2018 2508 2038 2511
rect 2050 2508 2054 2511
rect 2194 2508 2230 2511
rect 2386 2508 2406 2511
rect 2430 2508 2534 2511
rect 2538 2508 2542 2511
rect 2554 2508 2678 2511
rect 2770 2508 2806 2511
rect 2810 2508 2870 2511
rect 2882 2508 2886 2511
rect 3146 2508 3214 2511
rect 3226 2508 3310 2511
rect 3402 2508 3478 2511
rect 3634 2508 3670 2511
rect 3674 2508 3686 2511
rect 3690 2508 3718 2511
rect 3722 2508 3774 2511
rect 848 2503 850 2507
rect 854 2503 857 2507
rect 862 2503 864 2507
rect 1880 2503 1882 2507
rect 1886 2503 1889 2507
rect 1894 2503 1896 2507
rect 2430 2502 2433 2508
rect 2904 2503 2906 2507
rect 2910 2503 2913 2507
rect 2918 2503 2920 2507
rect 466 2498 630 2501
rect 1010 2498 1462 2501
rect 1466 2498 1590 2501
rect 1642 2498 1646 2501
rect 1674 2498 1678 2501
rect 1686 2498 1766 2501
rect 1930 2498 1958 2501
rect 1962 2498 2102 2501
rect 2106 2498 2150 2501
rect 2162 2498 2406 2501
rect 2426 2498 2430 2501
rect 2474 2498 2566 2501
rect 2570 2498 2598 2501
rect 2610 2498 2630 2501
rect 2730 2498 2894 2501
rect 3026 2498 3174 2501
rect 3178 2498 3638 2501
rect 934 2492 937 2498
rect 66 2488 366 2491
rect 386 2488 638 2491
rect 674 2488 926 2491
rect 942 2488 950 2491
rect 954 2488 998 2491
rect 1010 2488 1014 2491
rect 1122 2488 1206 2491
rect 1218 2488 1238 2491
rect 1398 2488 1406 2491
rect 1410 2488 1510 2491
rect 1522 2488 1526 2491
rect 1686 2491 1689 2498
rect 3654 2492 3657 2498
rect 1634 2488 1689 2491
rect 1818 2488 1862 2491
rect 1922 2488 1966 2491
rect 2242 2488 2286 2491
rect 2314 2488 2374 2491
rect 2426 2488 2582 2491
rect 2586 2488 2686 2491
rect 2794 2488 2814 2491
rect 2850 2488 2870 2491
rect 2898 2488 3118 2491
rect 3122 2488 3222 2491
rect 3242 2488 3246 2491
rect 3266 2488 3270 2491
rect 3306 2488 3326 2491
rect 3330 2488 3366 2491
rect 3386 2488 3438 2491
rect 3682 2488 3734 2491
rect 6 2481 9 2488
rect -26 2478 9 2481
rect 58 2478 102 2481
rect 242 2478 366 2481
rect 370 2478 486 2481
rect 602 2478 638 2481
rect 642 2478 710 2481
rect 810 2478 942 2481
rect 986 2478 1014 2481
rect 1094 2481 1097 2488
rect 1042 2478 1097 2481
rect 1170 2478 1206 2481
rect 1250 2478 1518 2481
rect 1522 2478 1686 2481
rect 1726 2481 1729 2488
rect 1698 2478 1729 2481
rect 1750 2481 1753 2488
rect 1750 2478 1830 2481
rect 1834 2478 1846 2481
rect 1898 2478 2006 2481
rect 2010 2478 2030 2481
rect 2206 2481 2209 2488
rect 2206 2478 2470 2481
rect 2486 2478 2494 2481
rect 2498 2478 2606 2481
rect 2614 2478 2622 2481
rect 2714 2478 2814 2481
rect 2826 2478 2841 2481
rect 2874 2478 2958 2481
rect 2982 2478 2990 2481
rect 2994 2478 3022 2481
rect 3090 2478 3134 2481
rect 3154 2478 3158 2481
rect 3162 2478 3198 2481
rect 3230 2481 3233 2488
rect 3230 2478 3246 2481
rect 3250 2478 3270 2481
rect 3294 2478 3366 2481
rect 3394 2478 3398 2481
rect 3522 2478 3542 2481
rect 3562 2478 3566 2481
rect 3586 2478 3590 2481
rect 3706 2478 3742 2481
rect -26 2472 -23 2478
rect -26 2468 -22 2472
rect 30 2471 33 2478
rect 10 2468 33 2471
rect 46 2468 86 2471
rect 378 2468 438 2471
rect 642 2468 678 2471
rect 690 2468 830 2471
rect 834 2468 897 2471
rect 930 2468 958 2471
rect 994 2468 998 2471
rect 1090 2468 1158 2471
rect 1402 2468 1438 2471
rect 1442 2468 1470 2471
rect 1506 2468 1558 2471
rect 1562 2468 1646 2471
rect 1730 2468 1758 2471
rect 1854 2471 1857 2478
rect 2614 2472 2617 2478
rect 2838 2472 2841 2478
rect 3062 2472 3065 2478
rect 3070 2472 3073 2478
rect 3294 2472 3297 2478
rect 1834 2468 1857 2471
rect 1962 2468 2078 2471
rect 2082 2468 2142 2471
rect 2146 2468 2198 2471
rect 2202 2468 2302 2471
rect 2630 2468 2694 2471
rect 2698 2468 2710 2471
rect 2738 2468 2750 2471
rect 2882 2468 2926 2471
rect 2986 2468 3006 2471
rect 3146 2468 3150 2471
rect 3250 2468 3270 2471
rect 3338 2468 3374 2471
rect 3386 2468 3390 2471
rect 3410 2468 3446 2471
rect 3482 2468 3486 2471
rect 3498 2468 3518 2471
rect 3694 2471 3697 2478
rect 3750 2472 3753 2478
rect 3694 2468 3750 2471
rect 22 2458 30 2461
rect 46 2461 49 2468
rect 190 2462 193 2468
rect 534 2462 537 2468
rect 34 2458 49 2461
rect 58 2458 62 2461
rect 442 2458 446 2461
rect 450 2458 473 2461
rect 686 2461 689 2468
rect 894 2462 897 2468
rect 686 2458 726 2461
rect 738 2458 742 2461
rect 770 2458 806 2461
rect 834 2458 838 2461
rect 906 2458 934 2461
rect 954 2458 958 2461
rect 970 2458 1030 2461
rect 1074 2458 1121 2461
rect 1138 2458 1150 2461
rect 1202 2458 1206 2461
rect 1314 2458 1406 2461
rect 1434 2458 1438 2461
rect 1514 2458 1534 2461
rect 1538 2458 1798 2461
rect 1842 2458 1894 2461
rect 1938 2458 1942 2461
rect 1954 2458 2062 2461
rect 2090 2458 2118 2461
rect 2226 2458 2350 2461
rect 2366 2461 2369 2468
rect 2366 2458 2390 2461
rect 2630 2461 2633 2468
rect 2450 2458 2633 2461
rect 2658 2458 2710 2461
rect 2746 2458 2750 2461
rect 2826 2458 2846 2461
rect 2850 2458 2854 2461
rect 2866 2458 2878 2461
rect 2906 2458 2950 2461
rect 2954 2458 2958 2461
rect 2978 2458 2998 2461
rect 3110 2461 3113 2468
rect 3110 2458 3414 2461
rect 3418 2458 3574 2461
rect 3614 2461 3617 2468
rect 3614 2458 3622 2461
rect 3650 2458 3702 2461
rect 470 2452 473 2458
rect 1118 2452 1121 2458
rect -26 2451 -22 2452
rect -26 2448 6 2451
rect 50 2448 65 2451
rect 90 2448 294 2451
rect 298 2448 454 2451
rect 474 2448 494 2451
rect 706 2448 718 2451
rect 722 2448 790 2451
rect 914 2448 934 2451
rect 1406 2451 1409 2458
rect 1854 2452 1857 2458
rect 1926 2452 1929 2458
rect 1210 2448 1233 2451
rect 1406 2448 1542 2451
rect 1546 2448 1710 2451
rect 1842 2448 1846 2451
rect 2042 2448 2081 2451
rect 62 2442 65 2448
rect 218 2438 438 2441
rect 602 2438 646 2441
rect 650 2438 782 2441
rect 870 2441 873 2448
rect 1230 2442 1233 2448
rect 2078 2442 2081 2448
rect 2182 2448 2206 2451
rect 2426 2448 2462 2451
rect 2482 2448 2694 2451
rect 2834 2448 2878 2451
rect 2986 2448 2990 2451
rect 2994 2448 3334 2451
rect 3346 2448 3350 2451
rect 3370 2448 3398 2451
rect 3402 2448 3470 2451
rect 3474 2448 3478 2451
rect 3506 2448 3534 2451
rect 3538 2448 3630 2451
rect 2182 2442 2185 2448
rect 786 2438 873 2441
rect 1058 2438 1110 2441
rect 1114 2438 1126 2441
rect 1130 2438 1134 2441
rect 1274 2438 1318 2441
rect 1322 2438 1534 2441
rect 1538 2438 1558 2441
rect 1570 2438 1702 2441
rect 2106 2438 2126 2441
rect 2290 2438 2310 2441
rect 2366 2441 2369 2448
rect 2366 2438 2438 2441
rect 2442 2438 2502 2441
rect 2706 2438 2798 2441
rect 2802 2438 3022 2441
rect 3058 2438 3134 2441
rect 3170 2438 3182 2441
rect 3186 2438 3214 2441
rect 3218 2438 3278 2441
rect 3330 2438 3438 2441
rect 3458 2438 3694 2441
rect 1422 2432 1425 2438
rect 314 2428 494 2431
rect 754 2428 838 2431
rect 914 2428 1182 2431
rect 1226 2428 1230 2431
rect 1546 2428 1566 2431
rect 1570 2428 1822 2431
rect 2126 2431 2129 2438
rect 2126 2428 2190 2431
rect 2250 2428 2302 2431
rect 2310 2431 2313 2438
rect 2310 2428 2718 2431
rect 2730 2428 2734 2431
rect 2786 2428 3062 2431
rect 3066 2428 3289 2431
rect 3362 2428 3414 2431
rect 3446 2431 3449 2438
rect 3446 2428 3510 2431
rect 178 2418 198 2421
rect 210 2418 790 2421
rect 1146 2418 1286 2421
rect 1290 2418 1494 2421
rect 1498 2418 1582 2421
rect 1586 2418 2022 2421
rect 2106 2418 2222 2421
rect 2282 2418 3070 2421
rect 3106 2418 3110 2421
rect 3130 2418 3166 2421
rect 3286 2421 3289 2428
rect 3622 2422 3625 2428
rect 3286 2418 3366 2421
rect 3670 2418 3678 2421
rect 3670 2412 3673 2418
rect 594 2408 654 2411
rect 1178 2408 1222 2411
rect 1282 2408 1334 2411
rect 1554 2408 1742 2411
rect 1810 2408 1814 2411
rect 1826 2408 2246 2411
rect 2266 2408 2358 2411
rect 2594 2408 3310 2411
rect 344 2403 346 2407
rect 350 2403 353 2407
rect 358 2403 360 2407
rect 1360 2403 1362 2407
rect 1366 2403 1369 2407
rect 1374 2403 1376 2407
rect 1470 2402 1473 2408
rect 2384 2403 2386 2407
rect 2390 2403 2393 2407
rect 2398 2403 2400 2407
rect 3408 2403 3410 2407
rect 3414 2403 3417 2407
rect 3422 2403 3424 2407
rect -26 2401 -22 2402
rect -26 2398 206 2401
rect 554 2398 942 2401
rect 946 2398 966 2401
rect 1018 2398 1254 2401
rect 1298 2398 1326 2401
rect 1482 2398 1745 2401
rect 1778 2398 1798 2401
rect 1802 2398 1950 2401
rect 1954 2398 2278 2401
rect 2438 2398 2470 2401
rect 2490 2398 2534 2401
rect 2730 2398 2814 2401
rect 2818 2398 2990 2401
rect 3082 2398 3294 2401
rect 3298 2398 3382 2401
rect 3626 2398 3742 2401
rect 558 2388 670 2391
rect 794 2388 910 2391
rect 1138 2388 1734 2391
rect 1742 2391 1745 2398
rect 1742 2388 1998 2391
rect 2042 2388 2166 2391
rect 2294 2388 2422 2391
rect 2438 2391 2441 2398
rect 2426 2388 2441 2391
rect 2778 2388 2830 2391
rect 2842 2388 2870 2391
rect 2994 2388 3262 2391
rect 3266 2388 3286 2391
rect 3466 2388 3526 2391
rect 3554 2388 3662 2391
rect 446 2381 449 2388
rect 558 2382 561 2388
rect 2294 2382 2297 2388
rect 446 2378 486 2381
rect 490 2378 494 2381
rect 618 2378 638 2381
rect 642 2378 758 2381
rect 898 2378 1030 2381
rect 1226 2378 1542 2381
rect 1578 2378 1590 2381
rect 1722 2378 1790 2381
rect 2522 2378 2558 2381
rect 2562 2378 2686 2381
rect 2690 2378 3206 2381
rect 3210 2378 3550 2381
rect 3602 2378 3614 2381
rect 3670 2381 3673 2388
rect 3670 2378 3702 2381
rect -26 2371 -22 2372
rect 30 2371 33 2378
rect -26 2368 33 2371
rect 526 2371 529 2378
rect 298 2368 529 2371
rect 546 2368 606 2371
rect 682 2368 686 2371
rect 778 2368 830 2371
rect 866 2368 950 2371
rect 1194 2368 2070 2371
rect 2074 2368 2510 2371
rect 2514 2368 2566 2371
rect 2618 2368 2758 2371
rect 2762 2368 2894 2371
rect 3026 2368 3030 2371
rect 3082 2368 3198 2371
rect 3218 2368 3230 2371
rect 3354 2368 3446 2371
rect 3482 2368 3558 2371
rect 3562 2368 3598 2371
rect 3666 2368 3710 2371
rect 3738 2368 3742 2371
rect 522 2358 622 2361
rect 670 2361 673 2368
rect 670 2358 718 2361
rect 834 2358 870 2361
rect 922 2358 926 2361
rect 950 2361 953 2368
rect 930 2358 1078 2361
rect 1274 2358 1310 2361
rect 1386 2358 1566 2361
rect 1602 2358 1606 2361
rect 1610 2358 1670 2361
rect 1698 2358 1702 2361
rect 1778 2358 1782 2361
rect 1794 2358 1814 2361
rect 1874 2358 1982 2361
rect 2026 2358 2030 2361
rect 2246 2358 2302 2361
rect 2362 2358 2550 2361
rect 2610 2358 2654 2361
rect 2658 2358 2665 2361
rect 2682 2358 2702 2361
rect 2738 2358 2958 2361
rect 3002 2358 3062 2361
rect 3066 2358 3078 2361
rect 3082 2358 3086 2361
rect 3090 2358 3118 2361
rect 3122 2358 3158 2361
rect 3162 2358 3302 2361
rect 3462 2361 3465 2368
rect 3450 2358 3694 2361
rect 3698 2358 3742 2361
rect 454 2352 457 2358
rect 742 2352 745 2358
rect -26 2351 -22 2352
rect -26 2348 6 2351
rect 218 2348 238 2351
rect 362 2348 382 2351
rect 458 2348 494 2351
rect 618 2348 646 2351
rect 666 2348 678 2351
rect 682 2348 694 2351
rect 762 2348 814 2351
rect 890 2348 894 2351
rect 994 2348 998 2351
rect 1074 2348 1118 2351
rect 1202 2348 1206 2351
rect 1210 2348 1366 2351
rect 1370 2348 1382 2351
rect 1386 2348 1414 2351
rect 1570 2348 1630 2351
rect 1634 2348 1662 2351
rect 1666 2348 1681 2351
rect 1690 2348 1774 2351
rect 1818 2348 1838 2351
rect 1842 2348 1846 2351
rect 1858 2348 1878 2351
rect 2246 2351 2249 2358
rect 2026 2348 2249 2351
rect 2258 2348 2286 2351
rect 2290 2348 2350 2351
rect 2490 2348 2574 2351
rect 2594 2348 2838 2351
rect 2882 2348 2894 2351
rect 3138 2348 3166 2351
rect 3210 2348 3214 2351
rect 3342 2351 3345 2358
rect 3342 2348 3382 2351
rect 3514 2348 3558 2351
rect 3602 2348 3686 2351
rect 3706 2348 3734 2351
rect 926 2342 929 2348
rect 450 2338 478 2341
rect 506 2338 510 2341
rect 514 2338 558 2341
rect 562 2338 702 2341
rect 722 2338 806 2341
rect 810 2338 878 2341
rect 938 2338 1230 2341
rect 1250 2338 1289 2341
rect 1298 2338 1310 2341
rect 1330 2338 1334 2341
rect 1578 2338 1670 2341
rect 1678 2341 1681 2348
rect 1678 2338 1694 2341
rect 1698 2338 1710 2341
rect 1806 2341 1809 2348
rect 1958 2342 1961 2348
rect 1786 2338 1809 2341
rect 1858 2338 1958 2341
rect 1966 2338 2014 2341
rect 2042 2338 2158 2341
rect 2314 2338 2321 2341
rect 2330 2338 2382 2341
rect 2422 2341 2425 2348
rect 2846 2342 2849 2348
rect 2854 2342 2857 2348
rect 2862 2342 2865 2348
rect 2998 2342 3001 2348
rect 3030 2342 3033 2348
rect 2418 2338 2425 2341
rect 2538 2338 2630 2341
rect 2666 2338 2702 2341
rect 2706 2338 2742 2341
rect 2754 2338 2798 2341
rect 2874 2338 2878 2341
rect 3066 2338 3118 2341
rect 3170 2338 3190 2341
rect 3250 2338 3278 2341
rect 3282 2338 3294 2341
rect 3458 2338 3550 2341
rect 3594 2338 3614 2341
rect 3634 2338 3742 2341
rect 430 2331 433 2338
rect 1286 2332 1289 2338
rect 430 2328 526 2331
rect 530 2328 678 2331
rect 690 2328 694 2331
rect 794 2328 1238 2331
rect 1266 2328 1270 2331
rect 1334 2328 1342 2331
rect 1382 2331 1385 2338
rect 1346 2328 1385 2331
rect 1478 2332 1481 2338
rect 1522 2328 1582 2331
rect 1618 2328 1638 2331
rect 1666 2328 1702 2331
rect 1818 2328 1846 2331
rect 1966 2331 1969 2338
rect 2438 2332 2441 2338
rect 2798 2332 2801 2338
rect 2806 2332 2809 2338
rect 1850 2328 1969 2331
rect 1994 2328 2046 2331
rect 2154 2328 2161 2331
rect 2338 2328 2342 2331
rect 2426 2328 2430 2331
rect 2482 2328 2590 2331
rect 2770 2328 2790 2331
rect 2982 2331 2985 2338
rect 3358 2332 3361 2338
rect 2834 2328 2985 2331
rect 3186 2328 3230 2331
rect 3250 2328 3270 2331
rect 3410 2328 3494 2331
rect 3498 2328 3542 2331
rect 3610 2328 3670 2331
rect 162 2318 870 2321
rect 906 2318 974 2321
rect 1050 2318 1190 2321
rect 1718 2321 1721 2328
rect 2158 2322 2161 2328
rect 1378 2318 1721 2321
rect 1726 2318 1870 2321
rect 1874 2318 1902 2321
rect 1922 2318 1982 2321
rect 2598 2321 2601 2328
rect 2178 2318 2601 2321
rect 2722 2318 2774 2321
rect 2830 2318 3038 2321
rect 3082 2318 3094 2321
rect 3098 2318 3158 2321
rect 3162 2318 3190 2321
rect 3226 2318 3342 2321
rect 3426 2318 3638 2321
rect 58 2308 62 2311
rect 66 2308 110 2311
rect 314 2308 326 2311
rect 370 2308 742 2311
rect 746 2308 806 2311
rect 810 2308 838 2311
rect 898 2308 926 2311
rect 1282 2308 1374 2311
rect 1726 2311 1729 2318
rect 1386 2308 1729 2311
rect 1738 2308 1846 2311
rect 1866 2308 1870 2311
rect 1946 2308 1974 2311
rect 2034 2308 2518 2311
rect 2830 2311 2833 2318
rect 2522 2308 2833 2311
rect 2930 2308 3006 2311
rect 3138 2308 3214 2311
rect 3546 2308 3582 2311
rect 3594 2308 3654 2311
rect 848 2303 850 2307
rect 854 2303 857 2307
rect 862 2303 864 2307
rect 1880 2303 1882 2307
rect 1886 2303 1889 2307
rect 1894 2303 1896 2307
rect 2904 2303 2906 2307
rect 2910 2303 2913 2307
rect 2918 2303 2920 2307
rect 466 2298 486 2301
rect 490 2298 550 2301
rect 738 2298 758 2301
rect 874 2298 1022 2301
rect 1098 2298 1390 2301
rect 1394 2298 1462 2301
rect 1594 2298 1873 2301
rect 2034 2298 2038 2301
rect 2066 2298 2582 2301
rect 2586 2298 2830 2301
rect 2850 2298 2862 2301
rect 3074 2298 3222 2301
rect 3234 2298 3342 2301
rect 3522 2298 3678 2301
rect 1018 2288 1105 2291
rect 1114 2288 1174 2291
rect 1226 2288 1406 2291
rect 1434 2288 1470 2291
rect 1502 2288 1758 2291
rect 1770 2288 1854 2291
rect 1870 2291 1873 2298
rect 1870 2288 1990 2291
rect 2002 2288 2046 2291
rect 2330 2288 2366 2291
rect 2378 2288 2422 2291
rect 2506 2288 2654 2291
rect 2658 2288 2734 2291
rect 2738 2288 2942 2291
rect 2950 2288 2958 2291
rect 2962 2288 2974 2291
rect 3050 2288 3230 2291
rect 3270 2288 3518 2291
rect 3566 2288 3574 2291
rect 3578 2288 3646 2291
rect 26 2278 30 2281
rect 326 2281 329 2288
rect 1102 2282 1105 2288
rect 202 2278 329 2281
rect 346 2278 462 2281
rect 1074 2278 1094 2281
rect 1114 2278 1118 2281
rect 1178 2278 1310 2281
rect 1414 2281 1417 2288
rect 1502 2282 1505 2288
rect 1734 2282 1737 2288
rect 2262 2282 2265 2288
rect 3270 2282 3273 2288
rect 3686 2282 3689 2288
rect 1414 2278 1502 2281
rect 1754 2278 1814 2281
rect 1866 2278 2118 2281
rect 2362 2278 2414 2281
rect 2426 2278 2462 2281
rect 2474 2278 2518 2281
rect 2650 2278 2846 2281
rect 2946 2278 3030 2281
rect 3042 2278 3110 2281
rect 3122 2278 3270 2281
rect 3282 2278 3286 2281
rect 3434 2278 3438 2281
rect 3458 2278 3462 2281
rect 3490 2278 3542 2281
rect 3570 2278 3574 2281
rect 18 2268 38 2271
rect 58 2268 102 2271
rect 114 2268 206 2271
rect 258 2268 414 2271
rect 682 2268 950 2271
rect 986 2268 1014 2271
rect 1018 2268 1246 2271
rect 1318 2271 1321 2278
rect 3734 2272 3737 2278
rect 1318 2268 1422 2271
rect 1450 2268 1454 2271
rect 1490 2268 1494 2271
rect 1506 2268 1518 2271
rect 1610 2268 1774 2271
rect 1794 2268 1798 2271
rect 1826 2268 1849 2271
rect 1866 2268 1870 2271
rect 1914 2268 1950 2271
rect 1954 2268 2006 2271
rect 2018 2268 2094 2271
rect 2098 2268 2126 2271
rect 2170 2268 2174 2271
rect 2378 2268 2382 2271
rect 2482 2268 2486 2271
rect 2498 2268 2558 2271
rect 2594 2268 2622 2271
rect 2634 2268 2638 2271
rect 2722 2268 2734 2271
rect 2778 2268 2822 2271
rect 2826 2268 2886 2271
rect 2890 2268 2950 2271
rect 3002 2268 3022 2271
rect 3042 2268 3046 2271
rect 3050 2268 3166 2271
rect 3202 2268 3206 2271
rect 3234 2268 3262 2271
rect 3370 2268 3398 2271
rect 3466 2268 3478 2271
rect 3538 2268 3710 2271
rect 98 2258 134 2261
rect 146 2258 150 2261
rect 202 2258 238 2261
rect 298 2258 390 2261
rect 482 2258 518 2261
rect 642 2258 694 2261
rect 826 2258 838 2261
rect 842 2258 862 2261
rect 890 2258 894 2261
rect 958 2261 961 2268
rect 958 2258 1006 2261
rect 1066 2258 1086 2261
rect 1114 2258 1126 2261
rect 1130 2258 1150 2261
rect 1154 2258 1294 2261
rect 1306 2258 1350 2261
rect 1370 2258 1382 2261
rect 1386 2258 1566 2261
rect 1570 2258 1582 2261
rect 1754 2258 1838 2261
rect 1846 2261 1849 2268
rect 2446 2262 2449 2268
rect 3334 2262 3337 2268
rect 1846 2258 1878 2261
rect 1882 2258 2118 2261
rect 2218 2258 2294 2261
rect 2298 2258 2358 2261
rect 2546 2258 2550 2261
rect 2586 2258 2614 2261
rect 2634 2258 2718 2261
rect 2786 2258 2846 2261
rect 2882 2258 2958 2261
rect 2986 2258 2990 2261
rect 3050 2258 3054 2261
rect 3106 2258 3118 2261
rect 3202 2258 3206 2261
rect 3274 2258 3294 2261
rect 3298 2258 3318 2261
rect 3386 2258 3454 2261
rect 3458 2258 3510 2261
rect 3526 2261 3529 2268
rect 3526 2258 3553 2261
rect 3586 2258 3606 2261
rect 3690 2258 3694 2261
rect 3730 2258 3766 2261
rect 1062 2252 1065 2258
rect 2614 2252 2617 2258
rect 3550 2252 3553 2258
rect -26 2251 -22 2252
rect -26 2248 6 2251
rect 26 2248 118 2251
rect 138 2248 246 2251
rect 914 2248 974 2251
rect 978 2248 1046 2251
rect 1074 2248 1078 2251
rect 1202 2248 1510 2251
rect 1530 2248 1550 2251
rect 1634 2248 1694 2251
rect 1730 2248 1750 2251
rect 1774 2248 1782 2251
rect 1842 2248 1846 2251
rect 1906 2248 1926 2251
rect 1930 2248 1998 2251
rect 2010 2248 2030 2251
rect 2090 2248 2102 2251
rect 2162 2248 2358 2251
rect 2410 2248 2486 2251
rect 2818 2248 2934 2251
rect 2986 2248 2998 2251
rect 3102 2248 3126 2251
rect 3138 2248 3166 2251
rect 3362 2248 3470 2251
rect 3474 2248 3478 2251
rect 3482 2248 3534 2251
rect 3562 2248 3566 2251
rect 3698 2248 3734 2251
rect 3754 2248 3761 2251
rect 1774 2242 1777 2248
rect 618 2238 638 2241
rect 1034 2238 1038 2241
rect 1042 2238 1134 2241
rect 1138 2238 1158 2241
rect 1210 2238 1246 2241
rect 1250 2238 1422 2241
rect 1530 2238 1758 2241
rect 1762 2238 1766 2241
rect 2046 2238 2278 2241
rect 2282 2238 2430 2241
rect 2442 2238 2470 2241
rect 2498 2238 2622 2241
rect 2934 2241 2937 2248
rect 3102 2242 3105 2248
rect 3758 2242 3761 2248
rect 2934 2238 3038 2241
rect 3330 2238 3374 2241
rect 3434 2238 3510 2241
rect 3554 2238 3574 2241
rect 3578 2238 3654 2241
rect 3658 2238 3662 2241
rect 3666 2238 3718 2241
rect 2022 2232 2025 2238
rect 2046 2232 2049 2238
rect 1138 2228 1142 2231
rect 1210 2228 1478 2231
rect 1482 2228 2006 2231
rect 2178 2228 3222 2231
rect 3250 2228 3326 2231
rect 3522 2228 3726 2231
rect 662 2221 665 2228
rect 290 2218 665 2221
rect 994 2218 1614 2221
rect 1818 2218 1958 2221
rect 2010 2218 2014 2221
rect 2018 2218 2326 2221
rect 2466 2218 2558 2221
rect 2626 2218 2822 2221
rect 2882 2218 3070 2221
rect 3226 2218 3494 2221
rect 3514 2218 3606 2221
rect 3646 2218 3654 2221
rect 3658 2218 3670 2221
rect 1974 2212 1977 2218
rect 90 2208 118 2211
rect 474 2208 590 2211
rect 762 2208 1166 2211
rect 1674 2208 1734 2211
rect 1746 2208 1814 2211
rect 2010 2208 2342 2211
rect 2346 2208 2350 2211
rect 2458 2208 2614 2211
rect 2618 2208 2910 2211
rect 2914 2208 3222 2211
rect 344 2203 346 2207
rect 350 2203 353 2207
rect 358 2203 360 2207
rect 1360 2203 1362 2207
rect 1366 2203 1369 2207
rect 1374 2203 1376 2207
rect 2384 2203 2386 2207
rect 2390 2203 2393 2207
rect 2398 2203 2400 2207
rect 3408 2203 3410 2207
rect 3414 2203 3417 2207
rect 3422 2203 3424 2207
rect 866 2198 990 2201
rect 1522 2198 1622 2201
rect 1626 2198 2150 2201
rect 2162 2198 2222 2201
rect 2250 2198 2374 2201
rect 2610 2198 3102 2201
rect 3106 2198 3398 2201
rect 34 2188 46 2191
rect 426 2188 630 2191
rect 826 2188 830 2191
rect 834 2188 1150 2191
rect 1226 2188 1230 2191
rect 1522 2188 1862 2191
rect 1930 2188 1966 2191
rect 1970 2188 1998 2191
rect 2002 2188 2174 2191
rect 2294 2188 2302 2191
rect 2306 2188 2318 2191
rect 2366 2188 2430 2191
rect 2462 2188 2518 2191
rect 2602 2188 2774 2191
rect 2778 2188 2806 2191
rect 2810 2188 2862 2191
rect 2906 2188 2998 2191
rect 3026 2188 3030 2191
rect 3338 2188 3406 2191
rect 3410 2188 3430 2191
rect 3458 2188 3494 2191
rect 3498 2188 3550 2191
rect 3554 2188 3590 2191
rect 3594 2188 3665 2191
rect 570 2178 574 2181
rect 602 2178 630 2181
rect 634 2178 662 2181
rect 666 2178 766 2181
rect 770 2178 838 2181
rect 1186 2178 1214 2181
rect 1218 2178 1342 2181
rect 1438 2181 1441 2188
rect 1438 2178 1502 2181
rect 1506 2178 1566 2181
rect 1570 2178 1686 2181
rect 1690 2178 1718 2181
rect 1770 2178 1790 2181
rect 1794 2178 2054 2181
rect 2162 2178 2222 2181
rect 2366 2181 2369 2188
rect 2278 2178 2369 2181
rect 2462 2182 2465 2188
rect 3662 2182 3665 2188
rect 2474 2178 2486 2181
rect 2642 2178 2662 2181
rect 2762 2178 2838 2181
rect 3090 2178 3198 2181
rect 3402 2178 3566 2181
rect 3586 2178 3598 2181
rect 550 2172 553 2178
rect 2278 2172 2281 2178
rect 554 2168 710 2171
rect 714 2168 774 2171
rect 778 2168 910 2171
rect 1106 2168 1126 2171
rect 1130 2168 1438 2171
rect 1650 2168 1766 2171
rect 2026 2168 2278 2171
rect 2378 2168 2462 2171
rect 2474 2168 2478 2171
rect 2514 2168 2814 2171
rect 3058 2168 3126 2171
rect 3250 2168 3270 2171
rect 3530 2168 3606 2171
rect 3610 2168 3710 2171
rect 526 2161 529 2168
rect 1558 2162 1561 2168
rect 1814 2162 1817 2168
rect 362 2158 529 2161
rect 546 2158 566 2161
rect 570 2158 590 2161
rect 594 2158 622 2161
rect 626 2158 721 2161
rect 738 2158 742 2161
rect 754 2158 758 2161
rect 802 2158 806 2161
rect 1106 2158 1110 2161
rect 1130 2158 1134 2161
rect 1450 2158 1470 2161
rect 1850 2158 1854 2161
rect 1918 2161 1921 2168
rect 1866 2158 1921 2161
rect 1950 2161 1953 2168
rect 1982 2162 1985 2168
rect 2294 2162 2297 2168
rect 1930 2158 1953 2161
rect 1962 2158 1966 2161
rect 2234 2158 2238 2161
rect 2434 2158 2462 2161
rect 2466 2158 2494 2161
rect 2506 2158 2510 2161
rect 2530 2158 2534 2161
rect 2674 2158 2678 2161
rect 2690 2158 2694 2161
rect 3114 2158 3126 2161
rect 3130 2158 3190 2161
rect 3194 2158 3214 2161
rect 3218 2158 3254 2161
rect 3258 2158 3302 2161
rect 3390 2161 3393 2168
rect 3606 2162 3609 2168
rect 3306 2158 3393 2161
rect 3418 2158 3430 2161
rect 3562 2158 3574 2161
rect 3682 2158 3686 2161
rect 3718 2161 3721 2168
rect 3698 2158 3721 2161
rect 718 2152 721 2158
rect -26 2151 -22 2152
rect -26 2148 6 2151
rect 426 2148 462 2151
rect 522 2148 526 2151
rect 634 2148 638 2151
rect 690 2148 710 2151
rect 722 2148 742 2151
rect 746 2148 798 2151
rect 802 2148 886 2151
rect 1018 2148 1198 2151
rect 1202 2148 1270 2151
rect 1466 2148 1470 2151
rect 1498 2148 1550 2151
rect 1618 2148 1670 2151
rect 1778 2148 1798 2151
rect 1802 2148 1902 2151
rect 1962 2148 1966 2151
rect 2182 2151 2185 2158
rect 1974 2148 2185 2151
rect 2210 2148 2614 2151
rect 2662 2151 2665 2158
rect 2658 2148 2665 2151
rect 2682 2148 2710 2151
rect 2746 2148 2782 2151
rect 2818 2148 2822 2151
rect 2850 2148 2862 2151
rect 2866 2148 2902 2151
rect 3110 2148 3150 2151
rect 3194 2148 3230 2151
rect 3266 2148 3294 2151
rect 3322 2148 3350 2151
rect 3482 2148 3502 2151
rect 3570 2148 3598 2151
rect 3618 2148 3638 2151
rect 3726 2151 3729 2158
rect 3714 2148 3729 2151
rect 134 2142 137 2148
rect 958 2142 961 2148
rect 1254 2142 1257 2148
rect 1310 2142 1313 2148
rect 1606 2142 1609 2148
rect 450 2138 454 2141
rect 530 2138 758 2141
rect 762 2138 822 2141
rect 826 2138 870 2141
rect 1042 2138 1046 2141
rect 1130 2138 1150 2141
rect 1178 2138 1190 2141
rect 1202 2138 1206 2141
rect 1418 2138 1454 2141
rect 1514 2138 1582 2141
rect 1618 2138 1638 2141
rect 1642 2138 1654 2141
rect 1666 2138 1798 2141
rect 1834 2138 1910 2141
rect 1974 2141 1977 2148
rect 2790 2142 2793 2148
rect 3110 2142 3113 2148
rect 1922 2138 1977 2141
rect 2250 2138 2310 2141
rect 2362 2138 2390 2141
rect 2434 2138 2446 2141
rect 2458 2138 2478 2141
rect 2530 2138 2718 2141
rect 2738 2138 2750 2141
rect 2754 2138 2785 2141
rect 2850 2138 2926 2141
rect 2962 2138 3038 2141
rect 3042 2138 3046 2141
rect 3082 2138 3086 2141
rect 3210 2138 3254 2141
rect 3314 2138 3393 2141
rect 3402 2138 3470 2141
rect 3626 2138 3734 2141
rect 118 2128 206 2131
rect 454 2131 457 2138
rect 2094 2132 2097 2138
rect 2206 2132 2209 2138
rect 2342 2132 2345 2138
rect 2782 2132 2785 2138
rect 370 2128 377 2131
rect 454 2128 502 2131
rect 594 2128 646 2131
rect 818 2128 1254 2131
rect 1294 2128 1310 2131
rect 1450 2128 1494 2131
rect 1498 2128 1518 2131
rect 1554 2128 1702 2131
rect 1706 2128 1886 2131
rect 1890 2128 1966 2131
rect 2226 2128 2254 2131
rect 2370 2128 2438 2131
rect 2450 2128 2470 2131
rect 2570 2128 2606 2131
rect 2730 2128 2769 2131
rect 2826 2128 2862 2131
rect 2882 2128 2886 2131
rect 2950 2131 2953 2138
rect 3158 2132 3161 2138
rect 2946 2128 2953 2131
rect 2962 2128 2966 2131
rect 3034 2128 3054 2131
rect 3066 2128 3086 2131
rect 3162 2128 3214 2131
rect 3218 2128 3310 2131
rect 3330 2128 3342 2131
rect 3390 2131 3393 2138
rect 3390 2128 3422 2131
rect 3530 2128 3534 2131
rect 3658 2128 3686 2131
rect 118 2122 121 2128
rect 374 2122 377 2128
rect 510 2121 513 2128
rect 1294 2122 1297 2128
rect 510 2118 566 2121
rect 938 2118 958 2121
rect 1394 2118 1446 2121
rect 1458 2118 1486 2121
rect 1702 2118 1750 2121
rect 1754 2118 1846 2121
rect 1874 2118 1878 2121
rect 1970 2118 2214 2121
rect 2446 2121 2449 2128
rect 2218 2118 2449 2121
rect 2518 2121 2521 2128
rect 2550 2122 2553 2128
rect 2766 2122 2769 2128
rect 2518 2118 2542 2121
rect 2594 2118 2686 2121
rect 2770 2118 2945 2121
rect 2954 2118 3046 2121
rect 3114 2118 3366 2121
rect 3650 2118 3678 2121
rect 3682 2118 3694 2121
rect 402 2108 758 2111
rect 762 2108 814 2111
rect 922 2108 942 2111
rect 1202 2108 1238 2111
rect 1274 2108 1278 2111
rect 1314 2108 1510 2111
rect 1522 2108 1558 2111
rect 1702 2111 1705 2118
rect 1586 2108 1705 2111
rect 1730 2108 1822 2111
rect 1826 2108 1862 2111
rect 1946 2108 2190 2111
rect 2194 2108 2422 2111
rect 2426 2108 2502 2111
rect 2506 2108 2526 2111
rect 2650 2108 2670 2111
rect 2738 2108 2894 2111
rect 2942 2111 2945 2118
rect 2942 2108 3022 2111
rect 3026 2108 3126 2111
rect 3226 2108 3230 2111
rect 3242 2108 3246 2111
rect 3322 2108 3342 2111
rect 3354 2108 3678 2111
rect 848 2103 850 2107
rect 854 2103 857 2107
rect 862 2103 864 2107
rect 1880 2103 1882 2107
rect 1886 2103 1889 2107
rect 1894 2103 1896 2107
rect 2904 2103 2906 2107
rect 2910 2103 2913 2107
rect 2918 2103 2920 2107
rect 3774 2102 3777 2108
rect 242 2098 262 2101
rect 442 2098 670 2101
rect 674 2098 718 2101
rect 1234 2098 1422 2101
rect 1498 2098 1614 2101
rect 1618 2098 1774 2101
rect 1786 2098 1870 2101
rect 1994 2098 2206 2101
rect 2274 2098 2334 2101
rect 2338 2098 2414 2101
rect 2418 2098 2481 2101
rect 2498 2098 2670 2101
rect 2698 2098 2734 2101
rect 2738 2098 2822 2101
rect 2930 2098 2990 2101
rect 3138 2098 3166 2101
rect 3170 2098 3198 2101
rect 3202 2098 3270 2101
rect 3274 2098 3334 2101
rect 3442 2098 3502 2101
rect 3682 2098 3726 2101
rect 506 2088 950 2091
rect 1138 2088 1182 2091
rect 1194 2088 1406 2091
rect 1426 2088 1534 2091
rect 1594 2088 1710 2091
rect 1770 2088 1926 2091
rect 1974 2091 1977 2098
rect 2478 2092 2481 2098
rect 1962 2088 1977 2091
rect 2002 2088 2222 2091
rect 2242 2088 2297 2091
rect 2306 2088 2350 2091
rect 2362 2088 2398 2091
rect 2418 2088 2430 2091
rect 2482 2088 2582 2091
rect 2586 2088 2598 2091
rect 2610 2088 2622 2091
rect 2666 2088 2734 2091
rect 2826 2088 2830 2091
rect 2854 2091 2857 2098
rect 2854 2088 2966 2091
rect 3130 2088 3606 2091
rect 3642 2088 3718 2091
rect 3746 2088 3750 2091
rect 398 2081 401 2088
rect 266 2078 401 2081
rect 450 2078 502 2081
rect 506 2078 654 2081
rect 890 2078 918 2081
rect 1130 2078 1134 2081
rect 1146 2078 1278 2081
rect 1406 2081 1409 2088
rect 2294 2082 2297 2088
rect 1406 2078 1462 2081
rect 1530 2078 1622 2081
rect 1626 2078 1641 2081
rect 1722 2078 1766 2081
rect 1810 2078 1830 2081
rect 1874 2078 1894 2081
rect 1914 2078 2070 2081
rect 2186 2078 2214 2081
rect 2306 2078 2310 2081
rect 2330 2078 2342 2081
rect 2350 2081 2353 2088
rect 2806 2082 2809 2088
rect 2350 2078 2406 2081
rect 2426 2078 2446 2081
rect 2450 2078 2526 2081
rect 2554 2078 2654 2081
rect 2730 2078 2782 2081
rect 2822 2081 2825 2088
rect 3094 2082 3097 2088
rect 2818 2078 2825 2081
rect 2834 2078 2950 2081
rect 2954 2078 3089 2081
rect 3162 2078 3190 2081
rect 3194 2078 3238 2081
rect 3306 2078 3334 2081
rect 3378 2078 3438 2081
rect 3458 2078 3462 2081
rect 3578 2078 3718 2081
rect 3766 2081 3769 2088
rect 3738 2078 3769 2081
rect -26 2071 -22 2072
rect 6 2071 9 2078
rect -26 2068 9 2071
rect 58 2068 78 2071
rect 222 2071 225 2078
rect 222 2068 230 2071
rect 274 2068 358 2071
rect 414 2071 417 2078
rect 414 2068 526 2071
rect 1030 2071 1033 2078
rect 810 2068 1033 2071
rect 1050 2068 1334 2071
rect 1338 2068 1358 2071
rect 1486 2071 1489 2078
rect 1638 2072 1641 2078
rect 1466 2068 1489 2071
rect 1746 2068 1790 2071
rect 1794 2068 1798 2071
rect 1802 2068 1862 2071
rect 1874 2068 1878 2071
rect 1890 2068 1934 2071
rect 2162 2068 2166 2071
rect 2226 2068 2454 2071
rect 2474 2068 2566 2071
rect 2578 2068 2582 2071
rect 2586 2068 2593 2071
rect 2602 2068 2662 2071
rect 2726 2071 2729 2078
rect 2674 2068 2729 2071
rect 2762 2068 2926 2071
rect 2994 2068 3054 2071
rect 3086 2071 3089 2078
rect 3086 2068 3246 2071
rect 3362 2068 3382 2071
rect 3386 2068 3446 2071
rect 3450 2068 3590 2071
rect 3594 2068 3630 2071
rect 66 2058 86 2061
rect 330 2058 486 2061
rect 746 2058 886 2061
rect 1154 2058 1214 2061
rect 1218 2058 1254 2061
rect 1446 2061 1449 2068
rect 1446 2058 1462 2061
rect 1502 2061 1505 2068
rect 1474 2058 1505 2061
rect 1582 2062 1585 2068
rect 1698 2058 1782 2061
rect 1802 2058 1825 2061
rect 1922 2058 1926 2061
rect 1978 2058 2222 2061
rect 2290 2058 2302 2061
rect 2314 2058 2446 2061
rect 2474 2058 2489 2061
rect 2546 2058 2566 2061
rect 2586 2058 2590 2061
rect 2618 2058 2694 2061
rect 2698 2058 2702 2061
rect 2778 2058 2942 2061
rect 2962 2058 3046 2061
rect 3106 2058 3110 2061
rect 3130 2058 3134 2061
rect 3294 2061 3297 2068
rect 3234 2058 3297 2061
rect 3302 2062 3305 2068
rect 3318 2062 3321 2068
rect 3362 2058 3390 2061
rect 3442 2058 3446 2061
rect 3546 2058 3566 2061
rect 3626 2058 3670 2061
rect 3742 2061 3745 2068
rect 3714 2058 3745 2061
rect 630 2052 633 2058
rect 1822 2052 1825 2058
rect 1942 2052 1945 2058
rect 2486 2052 2489 2058
rect 3046 2052 3049 2058
rect -26 2051 -22 2052
rect -26 2048 30 2051
rect 90 2048 318 2051
rect 474 2048 558 2051
rect 562 2048 598 2051
rect 802 2048 982 2051
rect 1146 2048 1177 2051
rect 1174 2042 1177 2048
rect 1394 2048 1454 2051
rect 1458 2048 1734 2051
rect 1770 2048 1782 2051
rect 1802 2048 1806 2051
rect 1866 2048 1902 2051
rect 2146 2048 2150 2051
rect 2178 2048 2182 2051
rect 2218 2048 2222 2051
rect 2354 2048 2486 2051
rect 2502 2048 2510 2051
rect 2514 2048 2590 2051
rect 2594 2048 2622 2051
rect 2666 2048 2697 2051
rect 2746 2048 2934 2051
rect 2978 2048 3030 2051
rect 3090 2048 3118 2051
rect 3242 2048 3262 2051
rect 3266 2048 3310 2051
rect 3362 2048 3374 2051
rect 3386 2048 3398 2051
rect 3474 2048 3542 2051
rect 3582 2051 3585 2058
rect 3570 2048 3670 2051
rect 3726 2048 3734 2051
rect 26 2038 97 2041
rect 458 2038 494 2041
rect 594 2038 678 2041
rect 906 2038 910 2041
rect 1206 2041 1209 2048
rect 1202 2038 1209 2041
rect 1218 2038 1470 2041
rect 1514 2038 1566 2041
rect 1742 2041 1745 2048
rect 2694 2042 2697 2048
rect 3726 2042 3729 2048
rect 1626 2038 1745 2041
rect 1778 2038 1830 2041
rect 1834 2038 2006 2041
rect 2114 2038 2382 2041
rect 2394 2038 2406 2041
rect 2442 2038 2470 2041
rect 2498 2038 2558 2041
rect 2602 2038 2662 2041
rect 2674 2038 2678 2041
rect 2898 2038 2990 2041
rect 2994 2038 3006 2041
rect 3018 2038 3038 2041
rect 3066 2038 3086 2041
rect 3130 2038 3478 2041
rect 3502 2038 3510 2041
rect 3514 2038 3526 2041
rect 3546 2038 3550 2041
rect 3642 2038 3646 2041
rect 3658 2038 3670 2041
rect 3738 2038 3742 2041
rect 94 2032 97 2038
rect 234 2028 590 2031
rect 602 2028 894 2031
rect 1174 2031 1177 2038
rect 1174 2028 1238 2031
rect 1554 2028 1750 2031
rect 1778 2028 1790 2031
rect 1858 2028 1926 2031
rect 1930 2028 1958 2031
rect 2430 2031 2433 2038
rect 1962 2028 2433 2031
rect 2482 2028 2894 2031
rect 2898 2028 3102 2031
rect 3370 2028 3374 2031
rect 3418 2028 3462 2031
rect 3466 2028 3526 2031
rect 3530 2028 3638 2031
rect 3690 2028 3745 2031
rect 138 2018 294 2021
rect 586 2018 694 2021
rect 738 2018 742 2021
rect 950 2012 953 2028
rect 3742 2022 3745 2028
rect 1162 2018 1294 2021
rect 1426 2018 1566 2021
rect 1810 2018 2622 2021
rect 2626 2018 2742 2021
rect 2810 2018 2830 2021
rect 2938 2018 2982 2021
rect 3010 2018 3190 2021
rect 3194 2018 3294 2021
rect 3314 2018 3486 2021
rect 3554 2018 3574 2021
rect 42 2008 270 2011
rect 530 2008 654 2011
rect 674 2008 694 2011
rect 714 2008 758 2011
rect 1018 2008 1174 2011
rect 1186 2008 1254 2011
rect 1442 2008 1654 2011
rect 1658 2008 1838 2011
rect 2146 2008 2278 2011
rect 2282 2008 2318 2011
rect 2330 2008 2374 2011
rect 2410 2008 2878 2011
rect 2882 2008 3214 2011
rect 3218 2008 3286 2011
rect 3490 2008 3526 2011
rect 3530 2008 3662 2011
rect 344 2003 346 2007
rect 350 2003 353 2007
rect 358 2003 360 2007
rect 1360 2003 1362 2007
rect 1366 2003 1369 2007
rect 1374 2003 1376 2007
rect 2384 2003 2386 2007
rect 2390 2003 2393 2007
rect 2398 2003 2400 2007
rect 3398 2002 3401 2008
rect 3408 2003 3410 2007
rect 3414 2003 3417 2007
rect 3422 2003 3424 2007
rect 162 1998 318 2001
rect 578 1998 598 2001
rect 778 1998 798 2001
rect 882 1998 950 2001
rect 1050 1998 1070 2001
rect 1162 1998 1182 2001
rect 1434 1998 1590 2001
rect 1594 1998 2230 2001
rect 2298 1998 2350 2001
rect 2354 1998 2374 2001
rect 2450 1998 2718 2001
rect 2746 1998 2998 2001
rect 3546 1998 3622 2001
rect 3642 1998 3758 2001
rect 1030 1992 1033 1998
rect -26 1991 -22 1992
rect -26 1988 14 1991
rect 514 1988 702 1991
rect 706 1988 886 1991
rect 1082 1988 1137 1991
rect 1134 1982 1137 1988
rect 1166 1988 1262 1991
rect 1266 1988 1318 1991
rect 1338 1988 1350 1991
rect 1418 1988 2022 1991
rect 2026 1988 2150 1991
rect 2250 1988 2398 1991
rect 2402 1988 2550 1991
rect 2554 1988 2838 1991
rect 2850 1988 2862 1991
rect 3146 1988 3222 1991
rect 3266 1988 3382 1991
rect 3394 1988 3614 1991
rect 1166 1982 1169 1988
rect 530 1978 574 1981
rect 1202 1978 1633 1981
rect -26 1971 -22 1972
rect 30 1971 33 1978
rect -26 1968 33 1971
rect 290 1968 358 1971
rect 362 1968 374 1971
rect 394 1968 566 1971
rect 642 1968 662 1971
rect 698 1968 934 1971
rect 962 1968 1057 1971
rect 1102 1971 1105 1978
rect 1074 1968 1126 1971
rect 1134 1971 1137 1978
rect 1630 1972 1633 1978
rect 1786 1978 1870 1981
rect 1874 1978 2030 1981
rect 2274 1978 2329 1981
rect 2370 1978 2510 1981
rect 2522 1978 2526 1981
rect 2570 1978 2598 1981
rect 2778 1978 3158 1981
rect 3162 1978 3646 1981
rect 1134 1968 1190 1971
rect 1218 1968 1230 1971
rect 1298 1968 1494 1971
rect 1758 1971 1761 1978
rect 2326 1972 2329 1978
rect 1746 1968 1761 1971
rect 1842 1968 1990 1971
rect 2362 1968 2430 1971
rect 2466 1968 2542 1971
rect 2642 1968 2694 1971
rect 2722 1968 2790 1971
rect 2874 1968 3294 1971
rect 3330 1968 3534 1971
rect 3594 1968 3606 1971
rect 3634 1968 3702 1971
rect 1054 1962 1057 1968
rect 26 1958 70 1961
rect 522 1958 609 1961
rect 618 1958 638 1961
rect 874 1958 910 1961
rect 994 1958 998 1961
rect 1058 1958 1110 1961
rect 1130 1958 1158 1961
rect 1202 1958 1310 1961
rect 1314 1958 1518 1961
rect 1582 1961 1585 1968
rect 1710 1962 1713 1968
rect 1582 1958 1606 1961
rect 1722 1958 1758 1961
rect 1818 1958 1830 1961
rect 1858 1958 2014 1961
rect 2026 1958 2190 1961
rect 2210 1958 2230 1961
rect 2266 1958 2270 1961
rect 2338 1958 2366 1961
rect 2410 1958 2438 1961
rect 2450 1958 2454 1961
rect 2522 1958 2574 1961
rect 2578 1958 2814 1961
rect 2866 1958 2894 1961
rect 2926 1958 2950 1961
rect 2954 1958 2961 1961
rect 2986 1958 3134 1961
rect 3154 1958 3174 1961
rect 3242 1958 3262 1961
rect 3394 1958 3398 1961
rect 3442 1958 3446 1961
rect 3514 1958 3518 1961
rect 3522 1958 3574 1961
rect 3578 1958 3590 1961
rect 3734 1961 3737 1968
rect 3674 1958 3737 1961
rect -26 1951 -22 1952
rect -26 1948 6 1951
rect 42 1948 49 1951
rect 46 1942 49 1948
rect 66 1948 70 1951
rect 74 1948 254 1951
rect 274 1948 558 1951
rect 606 1951 609 1958
rect 686 1952 689 1958
rect 2926 1952 2929 1958
rect 606 1948 630 1951
rect 642 1948 646 1951
rect 674 1948 681 1951
rect 722 1948 726 1951
rect 898 1948 982 1951
rect 994 1948 1078 1951
rect 1082 1948 1094 1951
rect 1098 1948 1142 1951
rect 1330 1948 1382 1951
rect 1474 1948 1478 1951
rect 1538 1948 1598 1951
rect 1610 1948 1662 1951
rect 1690 1948 1718 1951
rect 1826 1948 1830 1951
rect 1970 1948 1998 1951
rect 2234 1948 2270 1951
rect 2306 1948 2406 1951
rect 2410 1948 2414 1951
rect 2426 1948 2502 1951
rect 2506 1948 2590 1951
rect 2594 1948 2614 1951
rect 2634 1948 2710 1951
rect 2722 1948 2758 1951
rect 2762 1948 2766 1951
rect 2866 1948 2886 1951
rect 2954 1948 2974 1951
rect 3026 1948 3038 1951
rect 3050 1948 3054 1951
rect 3066 1948 3070 1951
rect 3078 1948 3150 1951
rect 3162 1948 3270 1951
rect 3310 1951 3313 1958
rect 3306 1948 3313 1951
rect 3330 1948 3334 1951
rect 3366 1948 3470 1951
rect 3478 1951 3481 1958
rect 3478 1948 3558 1951
rect 3562 1948 3606 1951
rect 3642 1948 3662 1951
rect 3666 1948 3670 1951
rect 54 1942 57 1948
rect 274 1938 310 1941
rect 314 1938 550 1941
rect 554 1938 566 1941
rect 586 1938 678 1941
rect 698 1938 742 1941
rect 922 1938 1014 1941
rect 1122 1938 1182 1941
rect 1186 1938 1222 1941
rect 1398 1941 1401 1948
rect 1846 1942 1849 1948
rect 1398 1938 1446 1941
rect 1570 1938 1590 1941
rect 1618 1938 1622 1941
rect 1634 1938 1638 1941
rect 1730 1938 1782 1941
rect 1866 1938 1974 1941
rect 1978 1938 1982 1941
rect 2126 1941 2129 1948
rect 2710 1942 2713 1948
rect 3078 1942 3081 1948
rect 3110 1942 3113 1948
rect 2126 1938 2198 1941
rect 2250 1938 2310 1941
rect 2330 1938 2350 1941
rect 2418 1938 2422 1941
rect 2434 1938 2446 1941
rect 2466 1938 2470 1941
rect 2482 1938 2526 1941
rect 2562 1938 2566 1941
rect 2602 1938 2606 1941
rect 2610 1938 2622 1941
rect 2658 1938 2702 1941
rect 2730 1938 2758 1941
rect 2762 1938 2798 1941
rect 2858 1938 2958 1941
rect 2962 1938 2974 1941
rect 3042 1938 3062 1941
rect 3154 1938 3158 1941
rect 3170 1938 3174 1941
rect 3282 1938 3286 1941
rect 3366 1941 3369 1948
rect 3306 1938 3369 1941
rect 3378 1938 3406 1941
rect 3466 1938 3486 1941
rect 3554 1938 3566 1941
rect 3610 1938 3654 1941
rect 3746 1938 3758 1941
rect 190 1932 193 1938
rect 2054 1932 2057 1938
rect 322 1928 465 1931
rect 482 1928 702 1931
rect 730 1928 742 1931
rect 754 1928 1014 1931
rect 1122 1928 1150 1931
rect 1154 1928 1174 1931
rect 1234 1928 1462 1931
rect 1514 1928 1526 1931
rect 1562 1928 1622 1931
rect 1626 1928 1718 1931
rect 1730 1928 1918 1931
rect 1922 1928 2030 1931
rect 2110 1931 2113 1938
rect 2110 1928 2126 1931
rect 2258 1928 2286 1931
rect 2322 1928 2446 1931
rect 2482 1928 2502 1931
rect 2506 1928 2686 1931
rect 2690 1928 2726 1931
rect 2730 1928 2750 1931
rect 2770 1928 2806 1931
rect 2882 1928 2894 1931
rect 2990 1931 2993 1938
rect 3446 1932 3449 1938
rect 2970 1928 2993 1931
rect 3002 1928 3086 1931
rect 3098 1928 3142 1931
rect 3194 1928 3246 1931
rect 3250 1928 3318 1931
rect 3322 1928 3326 1931
rect 3506 1928 3510 1931
rect 3530 1928 3558 1931
rect 3570 1928 3582 1931
rect 3634 1928 3662 1931
rect 462 1922 465 1928
rect 146 1918 174 1921
rect 178 1918 262 1921
rect 498 1918 622 1921
rect 818 1918 862 1921
rect 866 1918 902 1921
rect 954 1918 958 1921
rect 1322 1918 1390 1921
rect 1486 1918 1694 1921
rect 1722 1918 1774 1921
rect 2034 1918 2246 1921
rect 2258 1918 2422 1921
rect 2518 1918 2574 1921
rect 2698 1918 2710 1921
rect 2766 1921 2769 1928
rect 2738 1918 2769 1921
rect 2786 1918 2790 1921
rect 2794 1918 2838 1921
rect 2890 1918 2894 1921
rect 2906 1918 2958 1921
rect 2978 1918 3102 1921
rect 3142 1921 3145 1928
rect 3142 1918 3422 1921
rect 3426 1918 3446 1921
rect 774 1912 777 1918
rect 34 1908 110 1911
rect 114 1908 334 1911
rect 338 1908 446 1911
rect 466 1908 582 1911
rect 810 1908 838 1911
rect 946 1908 950 1911
rect 1486 1911 1489 1918
rect 2518 1912 2521 1918
rect 2966 1912 2969 1918
rect 1210 1908 1489 1911
rect 1562 1908 1582 1911
rect 1594 1908 1686 1911
rect 1698 1908 1790 1911
rect 1794 1908 1822 1911
rect 1938 1908 1950 1911
rect 1954 1908 1966 1911
rect 2106 1908 2118 1911
rect 2122 1908 2321 1911
rect 2330 1908 2366 1911
rect 2410 1908 2518 1911
rect 2538 1908 2814 1911
rect 2818 1908 2870 1911
rect 2938 1908 2950 1911
rect 3042 1908 3110 1911
rect 3130 1908 3166 1911
rect 3210 1908 3238 1911
rect 3258 1908 3262 1911
rect 3338 1908 3382 1911
rect 3418 1908 3454 1911
rect 848 1903 850 1907
rect 854 1903 857 1907
rect 862 1903 864 1907
rect 1880 1903 1882 1907
rect 1886 1903 1889 1907
rect 1894 1903 1896 1907
rect 98 1898 222 1901
rect 306 1898 494 1901
rect 498 1898 590 1901
rect 594 1898 790 1901
rect 906 1898 958 1901
rect 962 1898 1006 1901
rect 1394 1898 1526 1901
rect 1538 1898 1566 1901
rect 1578 1898 1646 1901
rect 1650 1898 1678 1901
rect 1682 1898 1750 1901
rect 1794 1898 1806 1901
rect 2298 1898 2310 1901
rect 2318 1901 2321 1908
rect 2904 1903 2906 1907
rect 2910 1903 2913 1907
rect 2918 1903 2920 1907
rect 2318 1898 2526 1901
rect 2730 1898 2782 1901
rect 2786 1898 2846 1901
rect 2850 1898 2862 1901
rect 2930 1898 3014 1901
rect 3042 1898 3046 1901
rect 3058 1898 3062 1901
rect 3090 1898 3158 1901
rect 3218 1898 3222 1901
rect 3234 1898 3254 1901
rect 3258 1898 3278 1901
rect 3290 1898 3310 1901
rect 3370 1898 3390 1901
rect 3450 1898 3662 1901
rect 470 1888 590 1891
rect 594 1888 958 1891
rect 1226 1888 1422 1891
rect 1490 1888 1526 1891
rect 1530 1888 1590 1891
rect 1602 1888 1622 1891
rect 1706 1888 1742 1891
rect 1746 1888 1870 1891
rect 2266 1888 2286 1891
rect 2294 1888 2430 1891
rect 2438 1888 2449 1891
rect 2474 1888 2686 1891
rect 2690 1888 2774 1891
rect 2794 1888 3049 1891
rect 3138 1888 3214 1891
rect 3222 1888 3246 1891
rect 3346 1888 3534 1891
rect 3570 1888 3590 1891
rect 3658 1888 3694 1891
rect 470 1882 473 1888
rect 130 1878 137 1881
rect 134 1872 137 1878
rect 370 1878 470 1881
rect 554 1878 558 1881
rect 570 1878 606 1881
rect 682 1878 694 1881
rect 706 1878 822 1881
rect 842 1878 929 1881
rect 938 1878 1062 1881
rect 1078 1881 1081 1888
rect 1066 1878 1081 1881
rect 1194 1878 1198 1881
rect 1214 1881 1217 1888
rect 1214 1878 1294 1881
rect 1306 1878 1414 1881
rect 1554 1878 1662 1881
rect 1674 1878 1726 1881
rect 1866 1878 1894 1881
rect 1954 1878 1966 1881
rect 2038 1881 2041 1888
rect 2294 1882 2297 1888
rect 2438 1882 2441 1888
rect 2446 1882 2449 1888
rect 3046 1882 3049 1888
rect 1974 1878 2041 1881
rect 2098 1878 2102 1881
rect 2274 1878 2278 1881
rect 2302 1878 2358 1881
rect 2362 1878 2422 1881
rect 2842 1878 2854 1881
rect 2858 1878 2881 1881
rect 2922 1878 2926 1881
rect 2962 1878 3038 1881
rect 3222 1881 3225 1888
rect 3114 1878 3225 1881
rect 3242 1878 3302 1881
rect 3306 1878 3310 1881
rect 3314 1878 3334 1881
rect 3386 1878 3422 1881
rect 3474 1878 3478 1881
rect 3506 1878 3574 1881
rect 3602 1878 3622 1881
rect 3642 1878 3686 1881
rect 3730 1878 3766 1881
rect 150 1871 153 1878
rect 926 1872 929 1878
rect 1510 1872 1513 1878
rect 150 1868 270 1871
rect 378 1868 510 1871
rect 514 1868 782 1871
rect 786 1868 918 1871
rect 962 1868 966 1871
rect 1002 1868 1054 1871
rect 1058 1868 1094 1871
rect 1146 1868 1190 1871
rect 1282 1868 1334 1871
rect 1522 1868 1526 1871
rect 1594 1868 1678 1871
rect 1806 1871 1809 1878
rect 1806 1868 1934 1871
rect 1974 1871 1977 1878
rect 2174 1872 2177 1878
rect 2302 1872 2305 1878
rect 2662 1872 2665 1878
rect 1962 1868 1977 1871
rect 2026 1868 2078 1871
rect 2202 1868 2294 1871
rect 2434 1868 2470 1871
rect 2506 1868 2550 1871
rect 2822 1871 2825 1878
rect 2794 1868 2825 1871
rect 2878 1872 2881 1878
rect 2986 1868 2998 1871
rect 3098 1868 3142 1871
rect 3154 1868 3166 1871
rect 3170 1868 3190 1871
rect 3194 1868 3278 1871
rect 3282 1868 3438 1871
rect 3482 1868 3486 1871
rect 3506 1868 3606 1871
rect 3642 1868 3654 1871
rect 3730 1868 3758 1871
rect 1334 1862 1337 1868
rect 2366 1862 2369 1868
rect 2942 1862 2945 1868
rect 210 1858 246 1861
rect 370 1858 406 1861
rect 458 1858 462 1861
rect 554 1858 590 1861
rect 634 1858 638 1861
rect 642 1858 726 1861
rect 746 1858 782 1861
rect 786 1858 790 1861
rect 898 1858 982 1861
rect 1034 1858 1070 1861
rect 1082 1858 1222 1861
rect 1226 1858 1238 1861
rect 1250 1858 1302 1861
rect 1434 1858 1438 1861
rect 1522 1858 2302 1861
rect 2306 1858 2342 1861
rect 2458 1858 2494 1861
rect 2522 1858 2526 1861
rect 2562 1858 2614 1861
rect 2770 1858 2774 1861
rect 2778 1858 2846 1861
rect 2874 1858 2878 1861
rect 2986 1858 3022 1861
rect 3122 1858 3238 1861
rect 3266 1858 3270 1861
rect 3338 1858 3342 1861
rect 3474 1858 3542 1861
rect 3694 1861 3697 1868
rect 3586 1858 3697 1861
rect -26 1851 -22 1852
rect -26 1848 6 1851
rect 306 1848 454 1851
rect 498 1848 598 1851
rect 618 1848 654 1851
rect 682 1848 718 1851
rect 770 1848 774 1851
rect 778 1848 790 1851
rect 858 1848 870 1851
rect 922 1848 958 1851
rect 1050 1848 1110 1851
rect 1186 1848 1438 1851
rect 1478 1851 1481 1858
rect 2414 1852 2417 1858
rect 3302 1852 3305 1858
rect 3374 1852 3377 1858
rect 3750 1852 3753 1858
rect 1478 1848 1614 1851
rect 1618 1848 1662 1851
rect 1666 1848 1686 1851
rect 1714 1848 1910 1851
rect 2018 1848 2070 1851
rect 2074 1848 2102 1851
rect 2234 1848 2310 1851
rect 2354 1848 2390 1851
rect 2530 1848 2606 1851
rect 2650 1848 2750 1851
rect 2770 1848 2798 1851
rect 2818 1848 2830 1851
rect 2938 1848 2942 1851
rect 2994 1848 3070 1851
rect 3162 1848 3174 1851
rect 3194 1848 3262 1851
rect 3498 1848 3510 1851
rect 3530 1848 3534 1851
rect 3594 1848 3630 1851
rect 1182 1842 1185 1848
rect 2454 1842 2457 1848
rect 466 1838 566 1841
rect 586 1838 814 1841
rect 906 1838 942 1841
rect 946 1838 990 1841
rect 994 1838 1182 1841
rect 1274 1838 1526 1841
rect 1538 1838 1566 1841
rect 1578 1838 1654 1841
rect 1954 1838 1958 1841
rect 1986 1838 2054 1841
rect 2058 1838 2262 1841
rect 2330 1838 2350 1841
rect 2354 1838 2406 1841
rect 2546 1838 2950 1841
rect 2994 1838 3086 1841
rect 3202 1838 3214 1841
rect 3258 1838 3278 1841
rect 3386 1838 3390 1841
rect 3526 1841 3529 1848
rect 3450 1838 3529 1841
rect 3558 1842 3561 1848
rect 3586 1838 3670 1841
rect 3698 1838 3710 1841
rect 3738 1838 3742 1841
rect 3762 1838 3822 1841
rect 490 1828 566 1831
rect 650 1828 654 1831
rect 706 1828 806 1831
rect 914 1828 998 1831
rect 1106 1828 1142 1831
rect 1146 1828 1150 1831
rect 1306 1828 1326 1831
rect 1330 1828 1582 1831
rect 1602 1828 1646 1831
rect 1650 1828 1894 1831
rect 1898 1828 2134 1831
rect 2570 1828 2958 1831
rect 2962 1828 3102 1831
rect 3122 1828 3150 1831
rect 3286 1831 3289 1838
rect 3226 1828 3289 1831
rect 3402 1828 3486 1831
rect 3546 1828 3614 1831
rect 3674 1828 3702 1831
rect 3706 1828 3758 1831
rect 410 1818 486 1821
rect 618 1818 734 1821
rect 810 1818 1158 1821
rect 1578 1818 1814 1821
rect 1818 1818 1990 1821
rect 1994 1818 2358 1821
rect 2378 1818 2486 1821
rect 2490 1818 2574 1821
rect 2578 1818 2766 1821
rect 2858 1818 3270 1821
rect 3394 1818 3718 1821
rect 530 1808 550 1811
rect 554 1808 582 1811
rect 946 1808 1078 1811
rect 1082 1808 1182 1811
rect 1554 1808 2150 1811
rect 2374 1811 2377 1818
rect 2226 1808 2377 1811
rect 2410 1808 2982 1811
rect 3010 1808 3022 1811
rect 3058 1808 3062 1811
rect 3066 1808 3078 1811
rect 3474 1808 3502 1811
rect 344 1803 346 1807
rect 350 1803 353 1807
rect 358 1803 360 1807
rect 1360 1803 1362 1807
rect 1366 1803 1369 1807
rect 1374 1803 1376 1807
rect 2384 1803 2386 1807
rect 2390 1803 2393 1807
rect 2398 1803 2400 1807
rect 3408 1803 3410 1807
rect 3414 1803 3417 1807
rect 3422 1803 3424 1807
rect 474 1798 630 1801
rect 826 1798 878 1801
rect 906 1798 1086 1801
rect 1554 1798 1574 1801
rect 1626 1798 1710 1801
rect 1834 1798 2006 1801
rect 2010 1798 2086 1801
rect 2554 1798 2678 1801
rect 2786 1798 2806 1801
rect 2826 1798 2838 1801
rect 2842 1798 3022 1801
rect 3242 1798 3318 1801
rect 3546 1798 3566 1801
rect 3594 1798 3742 1801
rect 2334 1792 2337 1798
rect 234 1788 686 1791
rect 690 1788 750 1791
rect 802 1788 974 1791
rect 1274 1788 1278 1791
rect 1290 1788 1601 1791
rect 1698 1788 1998 1791
rect 2002 1788 2126 1791
rect 2434 1788 2942 1791
rect 2946 1788 3238 1791
rect 3514 1788 3550 1791
rect 3602 1788 3774 1791
rect 1598 1782 1601 1788
rect 522 1778 574 1781
rect 722 1778 918 1781
rect 994 1778 1246 1781
rect 1458 1778 1582 1781
rect 1586 1778 1590 1781
rect 1610 1778 1670 1781
rect 1746 1778 1766 1781
rect 1786 1778 1798 1781
rect 1922 1778 2110 1781
rect 2114 1778 2278 1781
rect 2322 1778 3294 1781
rect 3298 1778 3654 1781
rect 330 1768 366 1771
rect 438 1771 441 1778
rect 438 1768 502 1771
rect 506 1768 526 1771
rect 570 1768 646 1771
rect 650 1768 686 1771
rect 698 1768 798 1771
rect 858 1768 982 1771
rect 1410 1768 1414 1771
rect 1418 1768 1454 1771
rect 1482 1768 1569 1771
rect 1642 1768 1910 1771
rect 1926 1768 1934 1771
rect 1938 1768 2030 1771
rect 2578 1768 2582 1771
rect 2650 1768 2702 1771
rect 2714 1768 2718 1771
rect 2762 1768 2886 1771
rect 2898 1768 2950 1771
rect 3122 1768 3166 1771
rect 3226 1768 3310 1771
rect 3354 1768 3382 1771
rect 3474 1768 3518 1771
rect 3530 1768 3606 1771
rect 3662 1771 3665 1778
rect 3662 1768 3670 1771
rect 1566 1762 1569 1768
rect 2118 1762 2121 1768
rect 2462 1762 2465 1768
rect 2510 1762 2513 1768
rect 3190 1762 3193 1768
rect 326 1758 358 1761
rect 450 1758 590 1761
rect 666 1758 758 1761
rect 802 1758 822 1761
rect 962 1758 998 1761
rect 1450 1758 1494 1761
rect 1610 1758 1625 1761
rect 1650 1758 1694 1761
rect 1794 1758 1798 1761
rect 1810 1758 1958 1761
rect 1962 1758 1974 1761
rect 2066 1758 2070 1761
rect 2194 1758 2230 1761
rect 2250 1758 2382 1761
rect 2530 1758 2638 1761
rect 2666 1758 2726 1761
rect 2778 1758 2854 1761
rect 2874 1758 2886 1761
rect 2922 1758 3030 1761
rect 3138 1758 3190 1761
rect 3306 1758 3358 1761
rect 3538 1758 3542 1761
rect 3562 1758 3590 1761
rect 3638 1761 3641 1768
rect 3610 1758 3646 1761
rect 3682 1758 3718 1761
rect 3742 1761 3745 1768
rect 3742 1758 3766 1761
rect 326 1752 329 1758
rect 790 1752 793 1758
rect -26 1751 -22 1752
rect -26 1748 6 1751
rect 194 1748 206 1751
rect 298 1748 302 1751
rect 306 1748 310 1751
rect 346 1748 382 1751
rect 466 1748 478 1751
rect 498 1748 534 1751
rect 546 1748 558 1751
rect 642 1748 657 1751
rect 674 1748 678 1751
rect 754 1748 769 1751
rect 818 1748 830 1751
rect 846 1751 849 1758
rect 846 1748 878 1751
rect 986 1748 1038 1751
rect 1374 1751 1377 1758
rect 1622 1752 1625 1758
rect 1234 1748 1382 1751
rect 1562 1748 1590 1751
rect 1594 1748 1606 1751
rect 1750 1751 1753 1758
rect 2862 1752 2865 1758
rect 3286 1752 3289 1758
rect 1730 1748 1838 1751
rect 1842 1748 1902 1751
rect 1906 1748 1950 1751
rect 1954 1748 1998 1751
rect 2090 1748 2542 1751
rect 2554 1748 2574 1751
rect 2626 1748 2630 1751
rect 2682 1748 2742 1751
rect 2762 1748 2798 1751
rect 2874 1748 2966 1751
rect 3074 1748 3078 1751
rect 3098 1748 3126 1751
rect 3162 1748 3166 1751
rect 3178 1748 3222 1751
rect 3226 1748 3233 1751
rect 3342 1748 3406 1751
rect 3434 1748 3446 1751
rect 3450 1748 3462 1751
rect 3490 1748 3518 1751
rect 3546 1748 3550 1751
rect 3570 1748 3630 1751
rect 3634 1748 3670 1751
rect 3698 1748 3734 1751
rect 3754 1748 3758 1751
rect 534 1742 537 1748
rect 654 1742 657 1748
rect 766 1742 769 1748
rect 2670 1742 2673 1748
rect 3342 1742 3345 1748
rect 314 1738 334 1741
rect 426 1738 462 1741
rect 666 1738 670 1741
rect 786 1738 806 1741
rect 922 1738 950 1741
rect 998 1738 1046 1741
rect 1050 1738 1054 1741
rect 1218 1738 1222 1741
rect 1498 1738 1566 1741
rect 1570 1738 1574 1741
rect 1586 1738 1622 1741
rect 1642 1738 1646 1741
rect 1658 1738 1830 1741
rect 1910 1738 1982 1741
rect 2026 1738 2070 1741
rect 2106 1738 2134 1741
rect 2162 1738 2294 1741
rect 2378 1738 2486 1741
rect 2522 1738 2526 1741
rect 2562 1738 2566 1741
rect 2586 1738 2657 1741
rect 2690 1738 2694 1741
rect 2706 1738 2710 1741
rect 2722 1738 2726 1741
rect 2786 1738 2790 1741
rect 2818 1738 2822 1741
rect 2882 1738 2942 1741
rect 2978 1738 2998 1741
rect 3250 1738 3294 1741
rect 3594 1738 3678 1741
rect 3698 1738 3702 1741
rect 134 1732 137 1738
rect 998 1732 1001 1738
rect 118 1728 126 1731
rect 290 1728 294 1731
rect 362 1728 374 1731
rect 378 1728 414 1731
rect 426 1728 430 1731
rect 434 1728 438 1731
rect 530 1728 662 1731
rect 682 1728 686 1731
rect 762 1728 774 1731
rect 794 1728 910 1731
rect 946 1728 950 1731
rect 1034 1728 1038 1731
rect 1066 1728 1094 1731
rect 1358 1731 1361 1738
rect 1162 1728 1361 1731
rect 1374 1732 1377 1738
rect 1622 1732 1625 1738
rect 1910 1732 1913 1738
rect 1982 1732 1985 1738
rect 2366 1732 2369 1738
rect 2550 1732 2553 1738
rect 1458 1728 1526 1731
rect 1698 1728 1750 1731
rect 1762 1728 1785 1731
rect 118 1722 121 1728
rect 1782 1722 1785 1728
rect 1842 1728 1902 1731
rect 1930 1728 1966 1731
rect 1994 1728 2022 1731
rect 2154 1728 2214 1731
rect 2218 1728 2286 1731
rect 2482 1728 2486 1731
rect 2578 1728 2638 1731
rect 2642 1728 2646 1731
rect 2654 1731 2657 1738
rect 2654 1728 2718 1731
rect 2746 1728 2990 1731
rect 3006 1731 3009 1738
rect 2994 1728 3009 1731
rect 3126 1732 3129 1738
rect 3146 1728 3278 1731
rect 3318 1731 3321 1738
rect 3282 1728 3321 1731
rect 3442 1728 3478 1731
rect 3690 1728 3694 1731
rect 490 1718 542 1721
rect 578 1718 622 1721
rect 626 1718 630 1721
rect 634 1718 694 1721
rect 754 1718 758 1721
rect 762 1718 830 1721
rect 834 1718 878 1721
rect 906 1718 926 1721
rect 938 1718 966 1721
rect 994 1718 1022 1721
rect 1034 1718 1038 1721
rect 1050 1718 1070 1721
rect 1178 1718 1318 1721
rect 1378 1718 1510 1721
rect 1814 1721 1817 1728
rect 1918 1722 1921 1728
rect 1814 1718 1854 1721
rect 2054 1721 2057 1728
rect 2054 1718 2126 1721
rect 2138 1718 2958 1721
rect 2970 1718 2974 1721
rect 2978 1718 3046 1721
rect 3058 1718 3062 1721
rect 3098 1718 3105 1721
rect 3210 1718 3374 1721
rect 3650 1718 3766 1721
rect 3102 1712 3105 1718
rect 274 1708 366 1711
rect 370 1708 486 1711
rect 738 1708 782 1711
rect 818 1708 830 1711
rect 882 1708 950 1711
rect 970 1708 1206 1711
rect 1242 1708 1486 1711
rect 1634 1708 1638 1711
rect 1778 1708 1870 1711
rect 1914 1708 1926 1711
rect 1930 1708 1942 1711
rect 1978 1708 2094 1711
rect 2106 1708 2398 1711
rect 2410 1708 2670 1711
rect 2674 1708 2686 1711
rect 2762 1708 2886 1711
rect 2954 1708 2974 1711
rect 2994 1708 3078 1711
rect 3226 1708 3254 1711
rect 3262 1708 3462 1711
rect 3546 1708 3574 1711
rect 3650 1708 3750 1711
rect 848 1703 850 1707
rect 854 1703 857 1707
rect 862 1703 864 1707
rect 1870 1702 1873 1708
rect 1880 1703 1882 1707
rect 1886 1703 1889 1707
rect 1894 1703 1896 1707
rect 2904 1703 2906 1707
rect 2910 1703 2913 1707
rect 2918 1703 2920 1707
rect 3262 1702 3265 1708
rect 450 1698 462 1701
rect 466 1698 494 1701
rect 498 1698 502 1701
rect 506 1698 598 1701
rect 602 1698 710 1701
rect 874 1698 1246 1701
rect 1266 1698 1377 1701
rect 1402 1698 1470 1701
rect 1522 1698 1606 1701
rect 1626 1698 1790 1701
rect 1810 1698 1838 1701
rect 1906 1698 1934 1701
rect 1938 1698 2054 1701
rect 2058 1698 2134 1701
rect 2146 1698 2198 1701
rect 2202 1698 2470 1701
rect 2474 1698 2598 1701
rect 2658 1698 2702 1701
rect 2770 1698 2798 1701
rect 2802 1698 2870 1701
rect 2962 1698 3206 1701
rect 3234 1698 3262 1701
rect 3330 1698 3630 1701
rect 3642 1698 3670 1701
rect 406 1691 409 1698
rect 394 1688 438 1691
rect 642 1688 745 1691
rect 770 1688 902 1691
rect 922 1688 942 1691
rect 1026 1688 1054 1691
rect 1066 1688 1070 1691
rect 1114 1688 1198 1691
rect 1234 1688 1238 1691
rect 1374 1691 1377 1698
rect 2710 1692 2713 1698
rect 1374 1688 1422 1691
rect 1482 1688 1529 1691
rect 1770 1688 1774 1691
rect 1842 1688 1894 1691
rect 1898 1688 1910 1691
rect 1986 1688 2030 1691
rect 2066 1688 2110 1691
rect 2370 1688 2374 1691
rect 2474 1688 2542 1691
rect 2554 1688 2678 1691
rect 2722 1688 2929 1691
rect 486 1681 489 1688
rect 742 1682 745 1688
rect 250 1678 377 1681
rect 486 1678 502 1681
rect 610 1678 662 1681
rect 778 1678 790 1681
rect 930 1678 934 1681
rect 1054 1681 1057 1688
rect 1526 1682 1529 1688
rect 938 1678 1118 1681
rect 1242 1678 1358 1681
rect 1466 1678 1518 1681
rect 1730 1678 1814 1681
rect 1858 1678 1870 1681
rect 1918 1681 1921 1688
rect 2230 1682 2233 1688
rect 1882 1678 1950 1681
rect 1954 1678 2022 1681
rect 2082 1678 2126 1681
rect 2298 1678 2310 1681
rect 2370 1678 2486 1681
rect 2594 1678 2646 1681
rect 2678 1681 2681 1688
rect 2926 1682 2929 1688
rect 3002 1688 3134 1691
rect 3162 1688 3246 1691
rect 3486 1688 3726 1691
rect 2650 1678 2657 1681
rect 2678 1678 2726 1681
rect 2730 1678 2742 1681
rect 2794 1678 2817 1681
rect 2850 1678 2854 1681
rect 2874 1678 2918 1681
rect 2982 1681 2985 1688
rect 3486 1682 3489 1688
rect 2982 1678 3006 1681
rect 3010 1678 3014 1681
rect 3050 1678 3070 1681
rect 3074 1678 3094 1681
rect 3106 1678 3142 1681
rect 3226 1678 3310 1681
rect 3314 1678 3334 1681
rect 3394 1678 3398 1681
rect 3530 1678 3542 1681
rect 3570 1678 3598 1681
rect 3650 1678 3678 1681
rect 94 1672 97 1678
rect -26 1671 -22 1672
rect -26 1668 6 1671
rect 218 1668 238 1671
rect 338 1668 366 1671
rect 374 1671 377 1678
rect 1182 1672 1185 1678
rect 1638 1672 1641 1678
rect 374 1668 622 1671
rect 650 1668 686 1671
rect 722 1668 742 1671
rect 834 1668 838 1671
rect 842 1668 1014 1671
rect 1030 1668 1038 1671
rect 1234 1668 1238 1671
rect 1322 1668 1334 1671
rect 1338 1668 1414 1671
rect 1434 1668 1470 1671
rect 1482 1668 1486 1671
rect 1506 1668 1510 1671
rect 1514 1668 1590 1671
rect 1682 1668 1726 1671
rect 1778 1668 1782 1671
rect 1850 1668 1918 1671
rect 1922 1668 1990 1671
rect 2010 1668 2038 1671
rect 2098 1668 2334 1671
rect 2338 1668 2406 1671
rect 2550 1671 2553 1678
rect 2814 1672 2817 1678
rect 2550 1668 2574 1671
rect 2642 1668 2662 1671
rect 2850 1668 2862 1671
rect 2914 1668 2974 1671
rect 2978 1668 2982 1671
rect 3002 1668 3166 1671
rect 3170 1668 3174 1671
rect 3234 1668 3238 1671
rect 3290 1668 3310 1671
rect 3322 1668 3326 1671
rect 3394 1668 3414 1671
rect 3418 1668 3518 1671
rect 3522 1668 3590 1671
rect 3594 1668 3670 1671
rect 3706 1668 3750 1671
rect 110 1662 113 1668
rect 1030 1662 1033 1668
rect 1110 1662 1113 1668
rect 170 1658 206 1661
rect 306 1658 334 1661
rect 338 1658 438 1661
rect 546 1658 598 1661
rect 666 1658 726 1661
rect 754 1658 766 1661
rect 802 1658 806 1661
rect 890 1658 902 1661
rect 938 1658 942 1661
rect 994 1658 998 1661
rect 1098 1658 1102 1661
rect 1210 1658 1342 1661
rect 1354 1658 1374 1661
rect 1386 1658 1566 1661
rect 1766 1661 1769 1668
rect 1674 1658 1769 1661
rect 1778 1658 1782 1661
rect 1810 1658 1814 1661
rect 1826 1658 1846 1661
rect 1890 1658 1918 1661
rect 2062 1661 2065 1668
rect 1962 1658 2065 1661
rect 2306 1658 2414 1661
rect 2490 1658 2582 1661
rect 2586 1658 2630 1661
rect 2650 1658 2686 1661
rect 2722 1658 2774 1661
rect 2778 1658 2782 1661
rect 2830 1661 2833 1668
rect 2826 1658 2833 1661
rect 3010 1658 3030 1661
rect 3366 1661 3369 1668
rect 3694 1662 3697 1668
rect 3138 1658 3430 1661
rect 3466 1658 3502 1661
rect 3506 1658 3510 1661
rect 3514 1658 3574 1661
rect 3578 1658 3646 1661
rect 3666 1658 3678 1661
rect 3722 1658 3734 1661
rect 3742 1658 3750 1661
rect 982 1652 985 1658
rect -26 1651 -22 1652
rect -26 1648 574 1651
rect 658 1648 678 1651
rect 682 1648 710 1651
rect 714 1648 734 1651
rect 754 1648 870 1651
rect 1002 1648 1006 1651
rect 1142 1651 1145 1658
rect 1142 1648 1454 1651
rect 1458 1648 1750 1651
rect 1754 1648 2118 1651
rect 2122 1648 2350 1651
rect 2378 1648 2566 1651
rect 2570 1648 2574 1651
rect 2674 1648 2734 1651
rect 2754 1648 2814 1651
rect 2826 1648 2838 1651
rect 3086 1651 3089 1658
rect 2874 1648 3049 1651
rect 3086 1648 3118 1651
rect 3162 1648 3166 1651
rect 3258 1648 3262 1651
rect 3394 1648 3526 1651
rect 3698 1648 3718 1651
rect 3742 1651 3745 1658
rect 3730 1648 3745 1651
rect 3754 1648 3758 1651
rect 3046 1642 3049 1648
rect 530 1638 686 1641
rect 690 1638 1158 1641
rect 1190 1638 1262 1641
rect 1314 1638 1334 1641
rect 1346 1638 1494 1641
rect 1786 1638 1862 1641
rect 1874 1638 1990 1641
rect 2114 1638 2662 1641
rect 2690 1638 3038 1641
rect 3182 1641 3185 1648
rect 3050 1638 3185 1641
rect 3234 1638 3238 1641
rect 3242 1638 3334 1641
rect 3338 1638 3358 1641
rect 3426 1638 3462 1641
rect 3490 1638 3534 1641
rect 3538 1638 3574 1641
rect 3674 1638 3734 1641
rect 3738 1638 3774 1641
rect 1190 1632 1193 1638
rect 354 1628 518 1631
rect 594 1628 606 1631
rect 610 1628 838 1631
rect 842 1628 1126 1631
rect 1130 1628 1174 1631
rect 1178 1628 1182 1631
rect 1262 1631 1265 1638
rect 1262 1628 1470 1631
rect 1474 1628 3502 1631
rect 3650 1628 3670 1631
rect 3746 1628 3758 1631
rect 514 1618 534 1621
rect 578 1618 1134 1621
rect 1166 1618 1174 1621
rect 1178 1618 1286 1621
rect 1290 1618 1302 1621
rect 1330 1618 1574 1621
rect 1762 1618 2358 1621
rect 2362 1618 2542 1621
rect 2610 1618 2710 1621
rect 2738 1618 3022 1621
rect 3026 1618 3302 1621
rect 3306 1618 3494 1621
rect 3562 1618 3710 1621
rect 602 1608 718 1611
rect 722 1608 750 1611
rect 762 1608 766 1611
rect 922 1608 1110 1611
rect 1234 1608 1254 1611
rect 1554 1608 1646 1611
rect 1658 1608 1846 1611
rect 1850 1608 1886 1611
rect 1930 1608 2286 1611
rect 2522 1608 2878 1611
rect 2994 1608 3054 1611
rect 3074 1608 3078 1611
rect 3090 1608 3198 1611
rect 344 1603 346 1607
rect 350 1603 353 1607
rect 358 1603 360 1607
rect 1350 1602 1353 1608
rect 1360 1603 1362 1607
rect 1366 1603 1369 1607
rect 1374 1603 1376 1607
rect 2384 1603 2386 1607
rect 2390 1603 2393 1607
rect 2398 1603 2400 1607
rect 3408 1603 3410 1607
rect 3414 1603 3417 1607
rect 3422 1603 3424 1607
rect 458 1598 614 1601
rect 618 1598 958 1601
rect 986 1598 998 1601
rect 1034 1598 1158 1601
rect 1234 1598 1238 1601
rect 1618 1598 1630 1601
rect 1666 1598 1958 1601
rect 1962 1598 2185 1601
rect 2194 1598 2366 1601
rect 2754 1598 2830 1601
rect 2890 1598 3070 1601
rect 3074 1598 3174 1601
rect 3490 1598 3494 1601
rect 3626 1598 3646 1601
rect 3650 1598 3702 1601
rect -26 1591 -22 1592
rect -26 1588 14 1591
rect 554 1588 697 1591
rect 730 1588 918 1591
rect 942 1588 950 1591
rect 954 1588 1270 1591
rect 1290 1588 1630 1591
rect 1634 1588 1734 1591
rect 1738 1588 2038 1591
rect 2042 1588 2094 1591
rect 2182 1591 2185 1598
rect 2182 1588 2646 1591
rect 3098 1588 3166 1591
rect 3170 1588 3214 1591
rect 3218 1588 3294 1591
rect 3298 1588 3454 1591
rect 3486 1588 3542 1591
rect 3642 1588 3734 1591
rect 470 1581 473 1588
rect 694 1582 697 1588
rect 1598 1582 1601 1588
rect 3486 1582 3489 1588
rect 194 1578 473 1581
rect 594 1578 670 1581
rect 754 1578 822 1581
rect 826 1578 1022 1581
rect 1154 1578 1222 1581
rect 1450 1578 1454 1581
rect 1466 1578 1486 1581
rect 1850 1578 1862 1581
rect 2162 1578 2662 1581
rect 2666 1578 2766 1581
rect 2946 1578 2998 1581
rect 3002 1578 3057 1581
rect 3114 1578 3134 1581
rect 3138 1578 3142 1581
rect 3190 1578 3366 1581
rect 3370 1578 3398 1581
rect 3450 1578 3478 1581
rect 3506 1578 3646 1581
rect -26 1571 -22 1572
rect 30 1571 33 1578
rect -26 1568 33 1571
rect 578 1568 646 1571
rect 670 1568 678 1571
rect 682 1568 694 1571
rect 722 1568 742 1571
rect 746 1568 870 1571
rect 986 1568 1166 1571
rect 1210 1568 1438 1571
rect 1442 1568 1518 1571
rect 1714 1568 2198 1571
rect 2202 1568 2230 1571
rect 2706 1568 2854 1571
rect 2894 1571 2897 1578
rect 2874 1568 2897 1571
rect 2922 1568 2982 1571
rect 3034 1568 3046 1571
rect 3054 1571 3057 1578
rect 3190 1572 3193 1578
rect 3054 1568 3110 1571
rect 3122 1568 3190 1571
rect 3226 1568 3310 1571
rect 3314 1568 3390 1571
rect 3394 1568 3422 1571
rect 3514 1568 3526 1571
rect 3546 1568 3574 1571
rect 3578 1568 3622 1571
rect 3738 1568 3758 1571
rect 298 1558 302 1561
rect 306 1558 318 1561
rect 382 1561 385 1568
rect 322 1558 385 1561
rect 442 1558 470 1561
rect 558 1561 561 1568
rect 498 1558 561 1561
rect 582 1558 686 1561
rect 898 1558 1046 1561
rect 1082 1558 1086 1561
rect 1194 1558 1406 1561
rect 1410 1558 1502 1561
rect 1770 1558 1873 1561
rect 1906 1558 2054 1561
rect 2058 1558 2350 1561
rect 2354 1558 2438 1561
rect 2442 1558 2454 1561
rect 2622 1561 2625 1568
rect 2594 1558 2625 1561
rect 2654 1561 2657 1568
rect 2654 1558 2734 1561
rect 2738 1558 2798 1561
rect 2818 1558 2846 1561
rect 2850 1558 2886 1561
rect 2890 1558 2942 1561
rect 3014 1561 3017 1568
rect 2970 1558 3017 1561
rect 3058 1558 3086 1561
rect 3122 1558 3126 1561
rect 3250 1558 3254 1561
rect 3258 1558 3278 1561
rect 3290 1558 3318 1561
rect 3498 1558 3534 1561
rect 3562 1558 3582 1561
rect 3614 1558 3654 1561
rect 3734 1561 3737 1568
rect 3730 1558 3737 1561
rect 582 1552 585 1558
rect -26 1551 -22 1552
rect -26 1548 6 1551
rect 346 1548 414 1551
rect 706 1548 734 1551
rect 826 1548 926 1551
rect 1054 1551 1057 1558
rect 1042 1548 1057 1551
rect 1466 1548 1558 1551
rect 1610 1548 1614 1551
rect 1634 1548 1742 1551
rect 1746 1548 1798 1551
rect 1870 1551 1873 1558
rect 1870 1548 1982 1551
rect 2098 1548 2102 1551
rect 2514 1548 2526 1551
rect 2602 1548 2630 1551
rect 2634 1548 2889 1551
rect 2898 1548 2910 1551
rect 3002 1548 3038 1551
rect 3078 1548 3086 1551
rect 3090 1548 3134 1551
rect 3154 1548 3222 1551
rect 3274 1548 3289 1551
rect 3358 1551 3361 1558
rect 3614 1552 3617 1558
rect 3354 1548 3361 1551
rect 3482 1548 3494 1551
rect 3514 1548 3518 1551
rect 3522 1548 3614 1551
rect 3658 1548 3678 1551
rect 3714 1548 3726 1551
rect 3730 1548 3742 1551
rect 462 1542 465 1548
rect 130 1538 158 1541
rect 330 1538 398 1541
rect 442 1538 454 1541
rect 466 1538 518 1541
rect 578 1538 590 1541
rect 610 1538 641 1541
rect 674 1538 878 1541
rect 890 1538 990 1541
rect 1114 1538 1198 1541
rect 1326 1541 1329 1548
rect 1326 1538 1382 1541
rect 1434 1538 1790 1541
rect 1802 1538 1830 1541
rect 2038 1541 2041 1548
rect 1970 1538 2041 1541
rect 2214 1541 2217 1548
rect 2130 1538 2217 1541
rect 2454 1541 2457 1548
rect 2454 1538 2550 1541
rect 2578 1538 2598 1541
rect 2834 1538 2870 1541
rect 2886 1541 2889 1548
rect 3286 1542 3289 1548
rect 2886 1538 2934 1541
rect 2986 1538 3078 1541
rect 3218 1538 3230 1541
rect 3234 1538 3238 1541
rect 3374 1541 3377 1548
rect 3354 1538 3377 1541
rect 3386 1538 3398 1541
rect 3470 1541 3473 1548
rect 3418 1538 3473 1541
rect 3530 1538 3606 1541
rect 3610 1538 3638 1541
rect 638 1532 641 1538
rect 298 1528 446 1531
rect 450 1528 462 1531
rect 714 1528 742 1531
rect 802 1528 806 1531
rect 830 1528 838 1531
rect 842 1528 902 1531
rect 954 1528 958 1531
rect 962 1528 974 1531
rect 1030 1531 1033 1538
rect 978 1528 1033 1531
rect 1058 1528 1190 1531
rect 1210 1528 1326 1531
rect 1498 1528 1545 1531
rect 1730 1528 1838 1531
rect 1866 1528 1870 1531
rect 1918 1531 1921 1538
rect 3310 1532 3313 1538
rect 1874 1528 1921 1531
rect 2250 1528 2278 1531
rect 2298 1528 2454 1531
rect 2506 1528 2526 1531
rect 2786 1528 2857 1531
rect 1446 1522 1449 1528
rect 1542 1522 1545 1528
rect 2022 1522 2025 1528
rect 2854 1522 2857 1528
rect 3042 1528 3102 1531
rect 3138 1528 3166 1531
rect 3170 1528 3238 1531
rect 3266 1528 3270 1531
rect 3322 1528 3486 1531
rect 3618 1528 3710 1531
rect 10 1518 494 1521
rect 498 1518 622 1521
rect 626 1518 750 1521
rect 754 1518 862 1521
rect 866 1518 894 1521
rect 898 1518 918 1521
rect 922 1518 926 1521
rect 1018 1518 1102 1521
rect 1114 1518 1326 1521
rect 1586 1518 1718 1521
rect 1734 1518 2017 1521
rect 2650 1518 2782 1521
rect 2974 1521 2977 1528
rect 3550 1522 3553 1528
rect 2874 1518 2977 1521
rect 3050 1518 3062 1521
rect 3066 1518 3222 1521
rect 3242 1518 3254 1521
rect 3306 1518 3342 1521
rect 3434 1518 3470 1521
rect 3626 1518 3638 1521
rect 66 1508 86 1511
rect 90 1508 262 1511
rect 386 1508 430 1511
rect 514 1508 718 1511
rect 730 1508 766 1511
rect 802 1508 830 1511
rect 882 1508 942 1511
rect 946 1508 1014 1511
rect 1146 1508 1174 1511
rect 1186 1508 1278 1511
rect 1290 1508 1342 1511
rect 1734 1511 1737 1518
rect 1530 1508 1737 1511
rect 2014 1511 2017 1518
rect 2014 1508 2150 1511
rect 2154 1508 2350 1511
rect 2714 1508 2734 1511
rect 2754 1508 2806 1511
rect 2810 1508 2814 1511
rect 2818 1508 2886 1511
rect 3074 1508 3230 1511
rect 3234 1508 3286 1511
rect 3298 1508 3302 1511
rect 3314 1508 3318 1511
rect 3338 1508 3342 1511
rect 3354 1508 3574 1511
rect 848 1503 850 1507
rect 854 1503 857 1507
rect 862 1503 864 1507
rect 1742 1502 1745 1508
rect 1880 1503 1882 1507
rect 1886 1503 1889 1507
rect 1894 1503 1896 1507
rect 2904 1503 2906 1507
rect 2910 1503 2913 1507
rect 2918 1503 2920 1507
rect 50 1498 302 1501
rect 410 1498 438 1501
rect 650 1498 726 1501
rect 970 1498 1150 1501
rect 1154 1498 1398 1501
rect 1458 1498 1502 1501
rect 1506 1498 1526 1501
rect 2250 1498 2366 1501
rect 2394 1498 2526 1501
rect 2746 1498 2846 1501
rect 2858 1498 2862 1501
rect 2926 1498 3094 1501
rect 3114 1498 3150 1501
rect 3158 1498 3182 1501
rect 3194 1498 3326 1501
rect 3330 1498 3494 1501
rect 3586 1498 3630 1501
rect 3634 1498 3670 1501
rect 162 1488 206 1491
rect 394 1488 462 1491
rect 530 1488 670 1491
rect 738 1488 790 1491
rect 842 1488 846 1491
rect 994 1488 1006 1491
rect 1090 1488 1094 1491
rect 1114 1488 1150 1491
rect 1170 1488 1174 1491
rect 1186 1488 1190 1491
rect 1354 1488 1358 1491
rect 1658 1488 1790 1491
rect 1810 1488 1838 1491
rect 1946 1488 1950 1491
rect 1970 1488 2174 1491
rect 2178 1488 2585 1491
rect 2602 1488 2609 1491
rect 2714 1488 2718 1491
rect 2926 1491 2929 1498
rect 2842 1488 2929 1491
rect 3026 1488 3030 1491
rect 3158 1491 3161 1498
rect 3034 1488 3161 1491
rect 3178 1488 3214 1491
rect 3218 1488 3398 1491
rect 3402 1488 3590 1491
rect 3618 1488 3702 1491
rect 262 1481 265 1488
rect 242 1478 265 1481
rect 382 1481 385 1488
rect 382 1478 390 1481
rect 402 1478 422 1481
rect 482 1478 513 1481
rect 522 1478 526 1481
rect 530 1478 534 1481
rect 630 1478 654 1481
rect 770 1478 966 1481
rect 994 1478 1006 1481
rect 1010 1478 1302 1481
rect 1306 1478 1310 1481
rect 1446 1481 1449 1488
rect 2582 1482 2585 1488
rect 2606 1482 2609 1488
rect 1346 1478 1902 1481
rect 1914 1478 2462 1481
rect 2466 1478 2574 1481
rect 2618 1478 2678 1481
rect 2682 1478 2750 1481
rect 2814 1481 2817 1488
rect 2762 1478 2817 1481
rect 2842 1478 3118 1481
rect 3162 1478 3166 1481
rect 3218 1478 3246 1481
rect 3266 1478 3454 1481
rect 3458 1478 3494 1481
rect 3538 1478 3542 1481
rect 3578 1478 3614 1481
rect 3658 1478 3678 1481
rect 3690 1478 3694 1481
rect 306 1468 414 1471
rect 426 1468 430 1471
rect 434 1468 486 1471
rect 510 1471 513 1478
rect 614 1471 617 1478
rect 510 1468 617 1471
rect 630 1472 633 1478
rect 2590 1472 2593 1478
rect 802 1468 814 1471
rect 842 1468 854 1471
rect 1050 1468 1054 1471
rect 1074 1468 1094 1471
rect 1146 1468 1198 1471
rect 1242 1468 1318 1471
rect 1370 1468 1537 1471
rect 1562 1468 1686 1471
rect 1706 1468 1766 1471
rect 1778 1468 1854 1471
rect 1858 1468 2094 1471
rect 2098 1468 2310 1471
rect 2338 1468 2366 1471
rect 2450 1468 2494 1471
rect 2602 1468 2606 1471
rect 2630 1470 2678 1471
rect -26 1458 753 1461
rect 802 1458 838 1461
rect 842 1458 934 1461
rect 938 1458 966 1461
rect 998 1461 1001 1468
rect 998 1458 1030 1461
rect 1058 1458 1062 1461
rect 1094 1461 1097 1468
rect 1206 1462 1209 1468
rect 1534 1462 1537 1468
rect 2246 1462 2249 1468
rect 1094 1458 1134 1461
rect 1138 1458 1150 1461
rect 1322 1458 1334 1461
rect 1554 1458 1558 1461
rect 1562 1458 1726 1461
rect 1730 1458 1758 1461
rect 1794 1458 1798 1461
rect 1810 1458 1870 1461
rect 1874 1458 1897 1461
rect 1906 1458 1910 1461
rect 2042 1458 2230 1461
rect 2330 1458 2398 1461
rect 2402 1458 2414 1461
rect 2418 1458 2470 1461
rect 2474 1458 2502 1461
rect 2510 1461 2513 1468
rect 2634 1468 2678 1470
rect 2682 1468 2846 1471
rect 2962 1468 2998 1471
rect 3018 1468 3062 1471
rect 3162 1468 3174 1471
rect 3218 1468 3294 1471
rect 3298 1468 3305 1471
rect 3370 1468 3462 1471
rect 3490 1468 3558 1471
rect 3650 1468 3662 1471
rect 3698 1468 3702 1471
rect 2510 1458 2566 1461
rect 2570 1458 2614 1461
rect 2730 1458 2942 1461
rect 2970 1458 2998 1461
rect 3002 1458 3006 1461
rect 3078 1458 3126 1461
rect 3130 1458 3158 1461
rect 3242 1458 3254 1461
rect 3266 1458 3454 1461
rect 3466 1458 3526 1461
rect 3530 1458 3534 1461
rect 3590 1461 3593 1468
rect 3550 1458 3593 1461
rect 3602 1458 3718 1461
rect 3762 1458 3774 1461
rect -26 1452 -23 1458
rect -26 1448 -22 1452
rect 18 1448 206 1451
rect 250 1448 406 1451
rect 430 1448 470 1451
rect 490 1448 494 1451
rect 594 1448 742 1451
rect 750 1451 753 1458
rect 750 1448 846 1451
rect 850 1448 953 1451
rect 1018 1448 1182 1451
rect 1210 1448 1270 1451
rect 1274 1448 1406 1451
rect 1450 1448 1550 1451
rect 1554 1448 1566 1451
rect 1634 1448 1638 1451
rect 1802 1448 1814 1451
rect 1882 1448 1886 1451
rect 1894 1451 1897 1458
rect 1934 1451 1937 1458
rect 3078 1452 3081 1458
rect 3550 1452 3553 1458
rect 1894 1448 1937 1451
rect 1946 1448 2038 1451
rect 2058 1448 2062 1451
rect 2306 1448 2310 1451
rect 2370 1448 2470 1451
rect 2474 1448 2478 1451
rect 2682 1448 2758 1451
rect 2762 1448 2798 1451
rect 2802 1448 2806 1451
rect 2954 1448 2982 1451
rect 3154 1448 3222 1451
rect 3362 1448 3374 1451
rect 3378 1448 3502 1451
rect 3562 1448 3622 1451
rect 3626 1448 3662 1451
rect 3698 1448 3758 1451
rect 3806 1451 3810 1452
rect 3778 1448 3810 1451
rect 430 1442 433 1448
rect 950 1442 953 1448
rect 458 1438 574 1441
rect 810 1438 822 1441
rect 1282 1438 1910 1441
rect 1914 1438 2078 1441
rect 2082 1438 2126 1441
rect 2426 1438 2446 1441
rect 2494 1441 2497 1448
rect 2494 1438 2534 1441
rect 2538 1438 2542 1441
rect 2610 1438 2654 1441
rect 2670 1441 2673 1448
rect 2670 1438 2686 1441
rect 2698 1438 3326 1441
rect 3330 1438 3622 1441
rect 3722 1438 3750 1441
rect 418 1428 446 1431
rect 450 1428 758 1431
rect 786 1428 814 1431
rect 854 1431 857 1438
rect 818 1428 857 1431
rect 958 1431 961 1438
rect 958 1428 1598 1431
rect 1602 1428 1838 1431
rect 2358 1431 2361 1438
rect 2358 1428 2486 1431
rect 2490 1428 2558 1431
rect 2722 1428 2798 1431
rect 2838 1428 3334 1431
rect 3338 1428 3446 1431
rect 3650 1428 3694 1431
rect 3698 1428 3745 1431
rect 170 1418 174 1421
rect 186 1418 726 1421
rect 754 1418 958 1421
rect 1082 1418 1086 1421
rect 1170 1418 1382 1421
rect 1466 1418 1566 1421
rect 1642 1418 1798 1421
rect 1802 1418 1822 1421
rect 1842 1418 2422 1421
rect 2838 1421 2841 1428
rect 3742 1422 3745 1428
rect 2434 1418 2841 1421
rect 2850 1418 2870 1421
rect 2874 1418 2894 1421
rect 3058 1418 3086 1421
rect 3130 1418 3198 1421
rect 3298 1418 3406 1421
rect 3714 1418 3726 1421
rect 74 1408 254 1411
rect 442 1408 518 1411
rect 802 1408 854 1411
rect 1450 1408 2358 1411
rect 2554 1408 2694 1411
rect 2802 1408 2846 1411
rect 2954 1408 3006 1411
rect 3018 1408 3038 1411
rect 3102 1408 3238 1411
rect 3634 1408 3734 1411
rect 344 1403 346 1407
rect 350 1403 353 1407
rect 358 1403 360 1407
rect 1360 1403 1362 1407
rect 1366 1403 1369 1407
rect 1374 1403 1376 1407
rect 2384 1403 2386 1407
rect 2390 1403 2393 1407
rect 2398 1403 2400 1407
rect 386 1398 550 1401
rect 570 1398 582 1401
rect 586 1398 598 1401
rect 754 1398 934 1401
rect 938 1398 942 1401
rect 1122 1398 1166 1401
rect 1226 1398 1350 1401
rect 1618 1398 1622 1401
rect 1794 1398 2070 1401
rect 2194 1398 2214 1401
rect 2226 1398 2230 1401
rect 2258 1398 2318 1401
rect 3102 1401 3105 1408
rect 3408 1403 3410 1407
rect 3414 1403 3417 1407
rect 3422 1403 3424 1407
rect 2562 1398 3105 1401
rect 3114 1398 3150 1401
rect 3154 1398 3286 1401
rect 3586 1398 3758 1401
rect 378 1388 510 1391
rect 666 1388 670 1391
rect 762 1388 806 1391
rect 810 1388 870 1391
rect 1314 1388 1382 1391
rect 1498 1388 1713 1391
rect 1722 1388 1878 1391
rect 1890 1388 2238 1391
rect 2362 1388 3046 1391
rect 3122 1388 3398 1391
rect 3402 1388 3486 1391
rect 3730 1388 3766 1391
rect -26 1381 -22 1382
rect 46 1381 49 1388
rect -26 1378 49 1381
rect 338 1378 646 1381
rect 730 1378 886 1381
rect 898 1378 1038 1381
rect 1178 1378 1446 1381
rect 1478 1381 1481 1388
rect 1710 1382 1713 1388
rect 1478 1378 1606 1381
rect 1770 1378 1918 1381
rect 1922 1378 2846 1381
rect 2890 1378 2894 1381
rect 2898 1378 3014 1381
rect 3118 1381 3121 1388
rect 3026 1378 3121 1381
rect 3130 1378 3134 1381
rect 3138 1378 3166 1381
rect 3330 1378 3566 1381
rect 3706 1378 3726 1381
rect 298 1368 382 1371
rect 498 1368 502 1371
rect 562 1368 582 1371
rect 682 1368 710 1371
rect 714 1368 790 1371
rect 794 1368 798 1371
rect 922 1368 1022 1371
rect 1170 1368 1486 1371
rect 1490 1368 1510 1371
rect 1646 1371 1649 1378
rect 1578 1368 1649 1371
rect 1742 1371 1745 1378
rect 1742 1368 1774 1371
rect 2010 1368 2121 1371
rect 2138 1368 2190 1371
rect 2194 1368 2270 1371
rect 2286 1368 2294 1371
rect 2298 1368 2382 1371
rect 2386 1368 2414 1371
rect 2418 1368 2510 1371
rect 2854 1371 2857 1378
rect 2794 1368 2857 1371
rect 2962 1368 2974 1371
rect 3018 1368 3110 1371
rect 3146 1368 3246 1371
rect 3258 1368 3342 1371
rect 3562 1368 3630 1371
rect 3634 1368 3742 1371
rect -26 1361 -22 1362
rect -26 1358 182 1361
rect 270 1361 273 1368
rect 1126 1362 1129 1368
rect 2118 1362 2121 1368
rect 270 1358 310 1361
rect 690 1358 710 1361
rect 714 1358 830 1361
rect 834 1358 838 1361
rect 946 1358 950 1361
rect 1418 1358 1438 1361
rect 1546 1358 1630 1361
rect 1634 1358 1662 1361
rect 1666 1358 1678 1361
rect 1754 1358 1766 1361
rect 1778 1358 1814 1361
rect 1818 1358 1878 1361
rect 2162 1358 2166 1361
rect 2274 1358 2286 1361
rect 2330 1358 2422 1361
rect 2498 1358 2502 1361
rect 2566 1361 2569 1368
rect 3774 1362 3777 1368
rect 2510 1358 2569 1361
rect 2762 1358 2766 1361
rect 2794 1358 2798 1361
rect 2874 1358 2878 1361
rect 2890 1358 2966 1361
rect 3002 1358 3022 1361
rect 3058 1358 3214 1361
rect 3218 1358 3294 1361
rect 3298 1358 3342 1361
rect 3346 1358 3390 1361
rect 3554 1358 3614 1361
rect 3674 1358 3766 1361
rect 258 1348 278 1351
rect 282 1348 302 1351
rect 474 1348 510 1351
rect 542 1351 545 1358
rect 1454 1352 1457 1358
rect 514 1348 545 1351
rect 602 1348 686 1351
rect 690 1348 758 1351
rect 826 1348 846 1351
rect 850 1348 910 1351
rect 914 1348 966 1351
rect 986 1348 990 1351
rect 1138 1348 1206 1351
rect 1274 1348 1406 1351
rect 1426 1348 1430 1351
rect 1502 1351 1505 1358
rect 2078 1352 2081 1358
rect 1474 1348 1505 1351
rect 1538 1348 1558 1351
rect 1562 1348 1638 1351
rect 1762 1348 1782 1351
rect 1834 1348 1846 1351
rect 2098 1348 2134 1351
rect 2138 1348 2190 1351
rect 2266 1348 2350 1351
rect 2354 1348 2438 1351
rect 2510 1351 2513 1358
rect 2466 1348 2513 1351
rect 2530 1348 2550 1351
rect 2562 1348 2582 1351
rect 2854 1351 2857 1358
rect 2818 1348 2857 1351
rect 2866 1348 2902 1351
rect 2906 1348 3006 1351
rect 3034 1348 3054 1351
rect 3058 1348 3065 1351
rect 3114 1348 3185 1351
rect 3202 1348 3206 1351
rect 3234 1348 3254 1351
rect 3338 1348 3345 1351
rect 3354 1348 3406 1351
rect 3510 1351 3513 1358
rect 3506 1348 3513 1351
rect 3578 1348 3598 1351
rect 3610 1348 3622 1351
rect 3650 1348 3654 1351
rect 3714 1348 3766 1351
rect 1070 1342 1073 1348
rect -26 1341 -22 1342
rect -26 1338 6 1341
rect 10 1338 30 1341
rect 530 1338 542 1341
rect 570 1338 590 1341
rect 594 1338 622 1341
rect 674 1338 774 1341
rect 778 1338 822 1341
rect 890 1338 934 1341
rect 954 1338 958 1341
rect 994 1338 1006 1341
rect 1246 1341 1249 1348
rect 1246 1338 1262 1341
rect 1702 1341 1705 1348
rect 3182 1342 3185 1348
rect 3318 1342 3321 1348
rect 3342 1342 3345 1348
rect 3446 1342 3449 1348
rect 3526 1342 3529 1348
rect 3542 1342 3545 1348
rect 1314 1338 1705 1341
rect 1738 1338 1841 1341
rect 1850 1338 2166 1341
rect 2170 1338 2198 1341
rect 2282 1338 2286 1341
rect 2330 1338 2358 1341
rect 2378 1338 2510 1341
rect 2514 1338 2574 1341
rect 2794 1338 2838 1341
rect 2866 1338 2870 1341
rect 2874 1338 3022 1341
rect 3026 1338 3062 1341
rect 3066 1338 3142 1341
rect 3370 1338 3374 1341
rect 3570 1338 3598 1341
rect 3606 1338 3614 1341
rect 3646 1338 3654 1341
rect 3658 1338 3694 1341
rect 174 1332 177 1338
rect 226 1328 334 1331
rect 546 1328 558 1331
rect 578 1328 686 1331
rect 834 1328 894 1331
rect 1018 1328 1089 1331
rect 1250 1328 1265 1331
rect 1354 1328 1366 1331
rect 1370 1328 1406 1331
rect 1442 1328 1526 1331
rect 1554 1328 1598 1331
rect 1618 1328 1622 1331
rect 1642 1328 1702 1331
rect 1722 1328 1734 1331
rect 1838 1331 1841 1338
rect 1838 1328 1862 1331
rect 1866 1328 2062 1331
rect 2130 1328 2134 1331
rect 2154 1328 2182 1331
rect 2210 1328 2238 1331
rect 2250 1328 2326 1331
rect 2330 1328 2406 1331
rect 2458 1328 2518 1331
rect 2546 1328 2574 1331
rect 2682 1328 2689 1331
rect 2874 1328 2942 1331
rect 2962 1328 2966 1331
rect 3018 1328 3030 1331
rect 3106 1328 3110 1331
rect 3114 1328 3222 1331
rect 3282 1328 3302 1331
rect 3306 1328 3358 1331
rect 3362 1328 3414 1331
rect 3482 1328 3582 1331
rect 3606 1331 3609 1338
rect 3598 1328 3609 1331
rect 3618 1328 3622 1331
rect 3650 1328 3750 1331
rect 1086 1322 1089 1328
rect 1262 1322 1265 1328
rect 2686 1322 2689 1328
rect 122 1318 398 1321
rect 402 1318 478 1321
rect 490 1318 542 1321
rect 698 1318 798 1321
rect 838 1318 918 1321
rect 930 1318 1006 1321
rect 1394 1318 1470 1321
rect 1522 1318 1534 1321
rect 1690 1318 1822 1321
rect 1914 1318 1926 1321
rect 1930 1318 2006 1321
rect 2042 1318 2254 1321
rect 2258 1318 2318 1321
rect 2322 1318 2398 1321
rect 2466 1318 2478 1321
rect 2530 1318 2534 1321
rect 2538 1318 2646 1321
rect 2842 1318 2990 1321
rect 3090 1318 3094 1321
rect 3138 1318 3142 1321
rect 3162 1318 3230 1321
rect 3234 1318 3358 1321
rect 3410 1318 3462 1321
rect 3466 1318 3486 1321
rect 3506 1318 3510 1321
rect 3518 1318 3526 1321
rect 3598 1321 3601 1328
rect 3530 1318 3601 1321
rect 3690 1318 3694 1321
rect 530 1308 534 1311
rect 838 1311 841 1318
rect 586 1308 841 1311
rect 890 1308 902 1311
rect 922 1308 966 1311
rect 1066 1308 1070 1311
rect 1090 1308 1094 1311
rect 1450 1308 1510 1311
rect 1562 1308 1726 1311
rect 1754 1308 1846 1311
rect 1906 1308 1934 1311
rect 2186 1308 2374 1311
rect 2402 1308 2478 1311
rect 2482 1308 2494 1311
rect 2646 1311 2649 1318
rect 2646 1308 2686 1311
rect 2802 1308 2886 1311
rect 2930 1308 2934 1311
rect 2970 1308 2998 1311
rect 3002 1308 3086 1311
rect 3178 1308 3222 1311
rect 3362 1308 3398 1311
rect 3418 1308 3454 1311
rect 3538 1308 3550 1311
rect 3586 1308 3670 1311
rect 848 1303 850 1307
rect 854 1303 857 1307
rect 862 1303 864 1307
rect 1880 1303 1882 1307
rect 1886 1303 1889 1307
rect 1894 1303 1896 1307
rect 2904 1303 2906 1307
rect 2910 1303 2913 1307
rect 2918 1303 2920 1307
rect 3174 1302 3177 1308
rect 450 1298 534 1301
rect 538 1298 590 1301
rect 674 1298 694 1301
rect 898 1298 990 1301
rect 1034 1298 1094 1301
rect 1106 1298 1142 1301
rect 1258 1298 1446 1301
rect 1474 1298 1566 1301
rect 1698 1298 1718 1301
rect 1834 1298 1838 1301
rect 2074 1298 2302 1301
rect 2306 1298 2334 1301
rect 2346 1298 2438 1301
rect 2458 1298 2646 1301
rect 2650 1298 2782 1301
rect 2786 1298 2814 1301
rect 2978 1298 2993 1301
rect 3010 1298 3105 1301
rect 3138 1298 3166 1301
rect 3194 1298 3230 1301
rect 3386 1298 3646 1301
rect 3682 1298 3726 1301
rect 2990 1292 2993 1298
rect 274 1288 438 1291
rect 466 1288 470 1291
rect 586 1288 734 1291
rect 786 1288 1030 1291
rect 1034 1288 1126 1291
rect 1402 1288 1641 1291
rect 1650 1288 1742 1291
rect 1810 1288 2086 1291
rect 2130 1288 2262 1291
rect 2274 1288 2286 1291
rect 2378 1288 2582 1291
rect 2826 1288 2830 1291
rect 2842 1288 2974 1291
rect 3074 1288 3094 1291
rect 3102 1291 3105 1298
rect 3190 1291 3193 1298
rect 3102 1288 3193 1291
rect 3290 1288 3350 1291
rect 3362 1288 3478 1291
rect 3546 1288 3582 1291
rect 3602 1288 3678 1291
rect 3690 1288 3758 1291
rect 402 1278 502 1281
rect 818 1278 926 1281
rect 962 1278 998 1281
rect 1142 1281 1145 1288
rect 1142 1278 1150 1281
rect 1362 1278 1406 1281
rect 1458 1278 1566 1281
rect 1638 1281 1641 1288
rect 2294 1282 2297 1288
rect 1638 1278 1854 1281
rect 1906 1278 1921 1281
rect 38 1272 41 1278
rect 382 1272 385 1278
rect 114 1268 158 1271
rect 162 1268 166 1271
rect 210 1268 342 1271
rect 482 1268 486 1271
rect 490 1268 518 1271
rect 702 1271 705 1278
rect 1390 1272 1393 1278
rect 1918 1272 1921 1278
rect 2354 1278 2398 1281
rect 2450 1278 2494 1281
rect 2498 1278 2542 1281
rect 2562 1278 2622 1281
rect 2626 1278 2630 1281
rect 2726 1281 2729 1288
rect 3214 1282 3217 1288
rect 2682 1278 2729 1281
rect 2834 1278 2950 1281
rect 2954 1278 2982 1281
rect 3066 1278 3110 1281
rect 3138 1278 3142 1281
rect 3242 1278 3310 1281
rect 3426 1278 3702 1281
rect 3722 1278 3742 1281
rect 702 1268 790 1271
rect 954 1268 1110 1271
rect 1154 1268 1158 1271
rect 1186 1268 1286 1271
rect 1530 1268 1606 1271
rect 1610 1268 1662 1271
rect 1698 1268 1702 1271
rect 1730 1268 1782 1271
rect 1786 1268 1846 1271
rect 1934 1271 1937 1278
rect 1934 1268 1942 1271
rect 1986 1268 2046 1271
rect 2234 1268 2238 1271
rect 2250 1268 2358 1271
rect 2362 1268 2374 1271
rect 2386 1268 2430 1271
rect 2434 1268 2486 1271
rect 2742 1271 2745 1278
rect 2742 1268 2774 1271
rect 2786 1268 2846 1271
rect 2850 1268 2902 1271
rect 3014 1271 3017 1278
rect 3342 1272 3345 1278
rect 3010 1268 3017 1271
rect 3050 1268 3134 1271
rect 3250 1268 3270 1271
rect 3282 1268 3318 1271
rect 3346 1268 3406 1271
rect 3418 1268 3422 1271
rect 3482 1268 3486 1271
rect 3514 1268 3582 1271
rect 3610 1268 3726 1271
rect 566 1261 569 1268
rect 1134 1262 1137 1268
rect 506 1258 569 1261
rect 746 1258 814 1261
rect 978 1258 1030 1261
rect 1082 1258 1086 1261
rect 1442 1258 1494 1261
rect 1502 1261 1505 1268
rect 1502 1258 1582 1261
rect 1586 1258 1718 1261
rect 1738 1258 2014 1261
rect 2050 1258 2086 1261
rect 2090 1258 2102 1261
rect 2250 1258 2270 1261
rect 2274 1258 2446 1261
rect 2522 1258 2526 1261
rect 2530 1258 2542 1261
rect 2574 1261 2577 1268
rect 2570 1258 2577 1261
rect 2618 1258 2622 1261
rect 2658 1258 2758 1261
rect 2762 1258 2846 1261
rect 2914 1258 2950 1261
rect 2970 1258 3062 1261
rect 3090 1258 3166 1261
rect 3170 1258 3246 1261
rect 3494 1261 3497 1268
rect 3378 1258 3497 1261
rect 3562 1258 3566 1261
rect 3634 1258 3638 1261
rect 3666 1258 3678 1261
rect 3690 1258 3726 1261
rect 3754 1258 3758 1261
rect 226 1248 302 1251
rect 778 1248 998 1251
rect 1002 1248 1198 1251
rect 1274 1248 1278 1251
rect 1406 1251 1409 1258
rect 3582 1252 3585 1258
rect 1406 1248 1526 1251
rect 1562 1248 1598 1251
rect 1650 1248 1750 1251
rect 1754 1248 1814 1251
rect 1858 1248 2534 1251
rect 2570 1248 2625 1251
rect 2650 1248 2878 1251
rect 2938 1248 2974 1251
rect 2978 1248 2982 1251
rect 3082 1248 3102 1251
rect 3146 1248 3230 1251
rect 3290 1248 3302 1251
rect 3394 1248 3446 1251
rect 3538 1248 3574 1251
rect 3602 1248 3734 1251
rect 2622 1242 2625 1248
rect 3750 1242 3753 1248
rect 170 1238 182 1241
rect 186 1238 206 1241
rect 266 1238 582 1241
rect 618 1238 774 1241
rect 1514 1238 1534 1241
rect 1738 1238 1758 1241
rect 1994 1238 1998 1241
rect 2170 1238 2302 1241
rect 2314 1238 2422 1241
rect 2626 1238 2841 1241
rect 2858 1238 3094 1241
rect 3098 1238 3206 1241
rect 3242 1238 3502 1241
rect 3506 1238 3574 1241
rect 3618 1238 3622 1241
rect 3690 1238 3694 1241
rect 626 1228 1110 1231
rect 1122 1228 1638 1231
rect 2614 1231 2617 1238
rect 2010 1228 2617 1231
rect 2838 1232 2841 1238
rect 3670 1232 3673 1238
rect 2994 1228 3334 1231
rect 3338 1228 3638 1231
rect 258 1218 374 1221
rect 458 1218 742 1221
rect 938 1218 1457 1221
rect 1466 1218 1518 1221
rect 1718 1221 1721 1228
rect 1650 1218 1721 1221
rect 1746 1218 2022 1221
rect 2026 1218 2038 1221
rect 2226 1218 2310 1221
rect 2322 1218 2622 1221
rect 3106 1218 3190 1221
rect 3426 1218 3617 1221
rect 3626 1218 3822 1221
rect 782 1208 1118 1211
rect 1454 1211 1457 1218
rect 1454 1208 1902 1211
rect 2242 1208 2294 1211
rect 2410 1208 2414 1211
rect 2458 1208 2494 1211
rect 2514 1208 2526 1211
rect 2530 1208 2958 1211
rect 2978 1208 3022 1211
rect 3082 1208 3182 1211
rect 3482 1208 3486 1211
rect 3614 1211 3617 1218
rect 3614 1208 3630 1211
rect 344 1203 346 1207
rect 350 1203 353 1207
rect 358 1203 360 1207
rect 90 1198 118 1201
rect 586 1198 638 1201
rect 782 1201 785 1208
rect 1360 1203 1362 1207
rect 1366 1203 1369 1207
rect 1374 1203 1376 1207
rect 2384 1203 2386 1207
rect 2390 1203 2393 1207
rect 2398 1203 2400 1207
rect 3408 1203 3410 1207
rect 3414 1203 3417 1207
rect 3422 1203 3424 1207
rect 642 1198 785 1201
rect 898 1198 1022 1201
rect 1026 1198 1134 1201
rect 1170 1198 1182 1201
rect 1186 1198 1353 1201
rect 1386 1198 1654 1201
rect 1658 1198 1686 1201
rect 1770 1198 2054 1201
rect 2642 1198 2646 1201
rect 2650 1198 2838 1201
rect 2842 1198 2942 1201
rect 2954 1198 2982 1201
rect 3170 1198 3182 1201
rect 3226 1198 3230 1201
rect 218 1188 254 1191
rect 890 1188 1270 1191
rect 1350 1191 1353 1198
rect 1766 1192 1769 1198
rect 3758 1192 3761 1198
rect 1350 1188 1478 1191
rect 1498 1188 1737 1191
rect 1930 1188 1934 1191
rect 1978 1188 2518 1191
rect 2522 1188 2742 1191
rect 2866 1188 2942 1191
rect 2946 1188 3062 1191
rect 3218 1188 3358 1191
rect 3366 1188 3510 1191
rect 686 1182 689 1188
rect 850 1178 886 1181
rect 1354 1178 1446 1181
rect 1522 1178 1662 1181
rect 1666 1178 1726 1181
rect 1734 1181 1737 1188
rect 1806 1182 1809 1188
rect 3366 1182 3369 1188
rect 1734 1178 1742 1181
rect 1746 1178 1774 1181
rect 1818 1178 1926 1181
rect 2258 1178 2334 1181
rect 2338 1178 2462 1181
rect 2466 1178 2854 1181
rect 2858 1178 2942 1181
rect 2946 1178 3270 1181
rect 3550 1181 3553 1188
rect 3550 1178 3606 1181
rect 430 1172 433 1178
rect -26 1171 -22 1172
rect -26 1168 6 1171
rect 234 1168 278 1171
rect 458 1168 478 1171
rect 482 1168 502 1171
rect 530 1168 542 1171
rect 570 1168 918 1171
rect 922 1168 1190 1171
rect 1330 1168 1390 1171
rect 1546 1168 1638 1171
rect 1738 1168 2142 1171
rect 2298 1168 2302 1171
rect 2426 1168 2462 1171
rect 2490 1168 2494 1171
rect 2594 1168 2606 1171
rect 2618 1168 2782 1171
rect 2810 1168 2822 1171
rect 2826 1168 2942 1171
rect 3066 1168 3126 1171
rect 3186 1168 3278 1171
rect 3494 1171 3497 1178
rect 3378 1168 3497 1171
rect 3546 1168 3550 1171
rect 3570 1168 3582 1171
rect 3726 1171 3729 1178
rect 3726 1168 3750 1171
rect 510 1162 513 1168
rect 2326 1162 2329 1168
rect 2950 1162 2953 1168
rect 74 1158 510 1161
rect 906 1158 1054 1161
rect 1194 1158 1414 1161
rect 1522 1158 1574 1161
rect 1626 1158 1774 1161
rect 1874 1158 1918 1161
rect 1922 1158 2142 1161
rect 2298 1158 2318 1161
rect 2354 1158 2358 1161
rect 2370 1158 2470 1161
rect 2474 1158 2478 1161
rect 2506 1158 2510 1161
rect 2554 1158 2598 1161
rect 2746 1158 2846 1161
rect 2866 1158 2902 1161
rect 2962 1158 2990 1161
rect 2994 1158 3030 1161
rect 3074 1158 3134 1161
rect 3162 1158 3198 1161
rect 3258 1158 3326 1161
rect 3330 1158 3342 1161
rect 3474 1158 3478 1161
rect 3586 1158 3614 1161
rect 3618 1158 3646 1161
rect 2150 1152 2153 1158
rect 3206 1152 3209 1158
rect -26 1151 -22 1152
rect -26 1148 6 1151
rect 186 1148 286 1151
rect 434 1148 438 1151
rect 458 1148 478 1151
rect 498 1148 542 1151
rect 546 1148 606 1151
rect 850 1148 862 1151
rect 874 1148 878 1151
rect 882 1148 910 1151
rect 930 1148 934 1151
rect 970 1148 990 1151
rect 1010 1148 1014 1151
rect 1082 1148 1126 1151
rect 1322 1148 1542 1151
rect 1546 1148 1558 1151
rect 1578 1148 1606 1151
rect 1626 1148 1678 1151
rect 1690 1148 1718 1151
rect 1722 1148 1750 1151
rect 1770 1148 1862 1151
rect 1866 1148 2033 1151
rect 2042 1148 2073 1151
rect 2306 1148 2310 1151
rect 2346 1148 2358 1151
rect 2378 1148 2430 1151
rect 2442 1148 2446 1151
rect 2466 1148 2630 1151
rect 2634 1148 2678 1151
rect 2786 1148 2870 1151
rect 2874 1148 2878 1151
rect 2962 1148 2966 1151
rect 2986 1148 3038 1151
rect 3042 1148 3118 1151
rect 3226 1148 3241 1151
rect 3322 1148 3366 1151
rect 3458 1148 3526 1151
rect 3530 1148 3534 1151
rect 3538 1148 3558 1151
rect 3562 1148 3742 1151
rect 1046 1142 1049 1148
rect 2030 1142 2033 1148
rect 2070 1142 2073 1148
rect 3238 1142 3241 1148
rect 70 1138 254 1141
rect 290 1138 342 1141
rect 438 1138 446 1141
rect 450 1138 537 1141
rect 70 1132 73 1138
rect 534 1132 537 1138
rect 810 1138 894 1141
rect 946 1138 990 1141
rect 994 1138 1022 1141
rect 1034 1138 1038 1141
rect 1082 1138 1086 1141
rect 1162 1138 1166 1141
rect 1258 1138 1326 1141
rect 1362 1138 1398 1141
rect 1402 1138 1470 1141
rect 1474 1138 1782 1141
rect 1798 1138 1814 1141
rect 1826 1138 1966 1141
rect 2322 1138 2374 1141
rect 2394 1138 2894 1141
rect 2902 1138 2998 1141
rect 3034 1138 3062 1141
rect 3074 1138 3158 1141
rect 3330 1138 3334 1141
rect 3338 1138 3350 1141
rect 3450 1138 3462 1141
rect 3482 1138 3614 1141
rect 3730 1138 3742 1141
rect 282 1128 313 1131
rect 550 1131 553 1138
rect 710 1132 713 1138
rect 550 1128 590 1131
rect 834 1128 942 1131
rect 1046 1131 1049 1138
rect 1246 1132 1249 1138
rect 1046 1128 1102 1131
rect 1342 1131 1345 1138
rect 1798 1132 1801 1138
rect 2214 1132 2217 1138
rect 1342 1128 1406 1131
rect 1410 1128 1414 1131
rect 1418 1128 1422 1131
rect 1434 1128 1438 1131
rect 1462 1128 1518 1131
rect 1530 1128 1534 1131
rect 1546 1128 1590 1131
rect 1594 1128 1614 1131
rect 1634 1128 1641 1131
rect 310 1122 313 1128
rect 346 1118 454 1121
rect 474 1118 478 1121
rect 482 1118 558 1121
rect 562 1118 710 1121
rect 1030 1121 1033 1128
rect 1262 1122 1265 1128
rect 1462 1122 1465 1128
rect 1638 1122 1641 1128
rect 1866 1128 1950 1131
rect 2026 1128 2209 1131
rect 2250 1128 2326 1131
rect 2330 1128 2358 1131
rect 2378 1128 2398 1131
rect 2434 1128 2457 1131
rect 2482 1128 2486 1131
rect 2514 1128 2542 1131
rect 2562 1128 2566 1131
rect 2578 1128 2606 1131
rect 2666 1128 2670 1131
rect 2754 1128 2814 1131
rect 2818 1128 2862 1131
rect 2902 1131 2905 1138
rect 2874 1128 2905 1131
rect 2970 1128 2990 1131
rect 2994 1128 2998 1131
rect 3010 1128 3038 1131
rect 3050 1128 3062 1131
rect 3166 1131 3169 1138
rect 3138 1128 3169 1131
rect 3190 1132 3193 1138
rect 3278 1132 3281 1138
rect 3234 1128 3246 1131
rect 3386 1128 3390 1131
rect 3426 1128 3454 1131
rect 3474 1128 3486 1131
rect 3634 1128 3646 1131
rect 762 1118 1025 1121
rect 1030 1118 1102 1121
rect 1162 1118 1246 1121
rect 1322 1118 1334 1121
rect 1338 1118 1382 1121
rect 1482 1118 1494 1121
rect 1546 1118 1574 1121
rect 1594 1118 1598 1121
rect 1610 1118 1630 1121
rect 1670 1121 1673 1128
rect 1670 1118 1854 1121
rect 1906 1118 2033 1121
rect 2042 1118 2046 1121
rect 2114 1118 2118 1121
rect 2162 1118 2174 1121
rect 2206 1121 2209 1128
rect 2454 1122 2457 1128
rect 2206 1118 2214 1121
rect 2314 1118 2342 1121
rect 2474 1118 2478 1121
rect 2494 1121 2497 1128
rect 2726 1122 2729 1128
rect 3126 1122 3129 1128
rect 3510 1122 3513 1128
rect 2490 1118 2497 1121
rect 2530 1118 2590 1121
rect 2594 1118 2598 1121
rect 2618 1118 2630 1121
rect 2642 1118 2662 1121
rect 2778 1118 2958 1121
rect 3010 1118 3030 1121
rect 3170 1118 3198 1121
rect 3202 1118 3214 1121
rect 3250 1118 3302 1121
rect 3426 1118 3430 1121
rect 3634 1118 3774 1121
rect 226 1108 262 1111
rect 266 1108 326 1111
rect 330 1108 422 1111
rect 426 1108 614 1111
rect 802 1108 830 1111
rect 1022 1111 1025 1118
rect 1022 1108 1238 1111
rect 1274 1108 1278 1111
rect 1482 1108 1870 1111
rect 1930 1108 1998 1111
rect 2030 1111 2033 1118
rect 2030 1108 2038 1111
rect 2042 1108 2166 1111
rect 2266 1108 2582 1111
rect 2586 1108 2598 1111
rect 2610 1108 2814 1111
rect 2946 1108 3022 1111
rect 3026 1108 3102 1111
rect 3106 1108 3110 1111
rect 3122 1108 3182 1111
rect 3494 1111 3497 1118
rect 3442 1108 3489 1111
rect 3494 1108 3518 1111
rect 3594 1108 3598 1111
rect 848 1103 850 1107
rect 854 1103 857 1107
rect 862 1103 864 1107
rect 1880 1103 1882 1107
rect 1886 1103 1889 1107
rect 1894 1103 1896 1107
rect 2904 1103 2906 1107
rect 2910 1103 2913 1107
rect 2918 1103 2920 1107
rect 2934 1102 2937 1108
rect 282 1098 318 1101
rect 322 1098 366 1101
rect 434 1098 462 1101
rect 746 1098 782 1101
rect 826 1098 838 1101
rect 970 1098 1022 1101
rect 1090 1098 1166 1101
rect 1170 1098 1206 1101
rect 1210 1098 1830 1101
rect 1946 1098 2286 1101
rect 2290 1098 2742 1101
rect 3026 1098 3230 1101
rect 3486 1101 3489 1108
rect 3486 1098 3542 1101
rect 3650 1098 3686 1101
rect 3462 1092 3465 1098
rect 242 1088 310 1091
rect 338 1088 454 1091
rect 698 1088 822 1091
rect 842 1088 974 1091
rect 986 1088 1566 1091
rect 1570 1088 1678 1091
rect 1682 1088 1710 1091
rect 2002 1088 2081 1091
rect 2090 1088 2110 1091
rect 2130 1088 2305 1091
rect 134 1081 137 1088
rect 134 1078 158 1081
rect 194 1078 230 1081
rect 614 1081 617 1088
rect 242 1078 617 1081
rect 714 1078 974 1081
rect 998 1078 1030 1081
rect 1122 1078 1126 1081
rect 1154 1078 1158 1081
rect 1218 1078 1222 1081
rect 1234 1078 1238 1081
rect 1266 1078 1318 1081
rect 1466 1078 1494 1081
rect 1626 1078 1662 1081
rect 1674 1078 1678 1081
rect 1682 1078 1766 1081
rect 1774 1081 1777 1088
rect 1774 1078 1878 1081
rect 1894 1081 1897 1088
rect 1894 1078 1902 1081
rect 1962 1078 2054 1081
rect 2078 1081 2081 1088
rect 2302 1082 2305 1088
rect 2346 1088 2446 1091
rect 2458 1088 2558 1091
rect 2646 1088 2654 1091
rect 2658 1088 2670 1091
rect 2682 1088 2694 1091
rect 2698 1088 2750 1091
rect 2762 1088 2782 1091
rect 2946 1088 3014 1091
rect 3038 1088 3094 1091
rect 3122 1088 3190 1091
rect 3330 1088 3334 1091
rect 3590 1088 3598 1091
rect 3602 1088 3686 1091
rect 2326 1082 2329 1088
rect 2078 1078 2086 1081
rect 2090 1078 2094 1081
rect 2202 1078 2206 1081
rect 2354 1078 2406 1081
rect 2418 1078 2494 1081
rect 2498 1078 2502 1081
rect 2598 1081 2601 1088
rect 2522 1078 2601 1081
rect 2610 1078 2638 1081
rect 2642 1078 2646 1081
rect 2650 1078 2710 1081
rect 2714 1078 2830 1081
rect 3038 1081 3041 1088
rect 3246 1082 3249 1088
rect 2866 1078 3041 1081
rect 3082 1078 3142 1081
rect 3146 1078 3190 1081
rect 3250 1078 3470 1081
rect 3474 1078 3502 1081
rect 3530 1078 3550 1081
rect 3570 1078 3590 1081
rect 3706 1078 3734 1081
rect -26 1071 -22 1072
rect 30 1071 33 1078
rect -26 1068 33 1071
rect 158 1071 161 1078
rect 998 1072 1001 1078
rect 158 1068 438 1071
rect 554 1068 694 1071
rect 826 1068 886 1071
rect 906 1068 958 1071
rect 978 1068 985 1071
rect 1102 1071 1105 1078
rect 1342 1072 1345 1078
rect 1558 1072 1561 1078
rect 1102 1068 1334 1071
rect 1450 1068 1558 1071
rect 1594 1068 1638 1071
rect 1650 1068 1790 1071
rect 1938 1068 1998 1071
rect 2074 1068 2174 1071
rect 2178 1068 2182 1071
rect 2194 1068 2230 1071
rect 2370 1068 2430 1071
rect 2482 1068 2526 1071
rect 2546 1068 2598 1071
rect 2610 1068 2657 1071
rect 2674 1068 2686 1071
rect 2722 1068 2758 1071
rect 2762 1068 2814 1071
rect 2838 1071 2841 1078
rect 3606 1072 3609 1078
rect 2838 1068 2854 1071
rect 2858 1068 2862 1071
rect 2978 1068 3150 1071
rect 3226 1068 3286 1071
rect 3290 1068 3342 1071
rect 3354 1068 3358 1071
rect 3426 1068 3430 1071
rect 3466 1068 3486 1071
rect 3506 1068 3534 1071
rect 3682 1068 3710 1071
rect 3714 1068 3774 1071
rect 982 1062 985 1068
rect 26 1058 30 1061
rect 50 1058 54 1061
rect 234 1058 246 1061
rect 250 1058 294 1061
rect 302 1058 318 1061
rect 338 1058 718 1061
rect 754 1058 774 1061
rect 938 1058 942 1061
rect 1014 1061 1017 1068
rect 1002 1058 1017 1061
rect 1034 1058 1110 1061
rect 1146 1058 1262 1061
rect 1418 1058 1470 1061
rect 1482 1058 1502 1061
rect 1506 1058 1510 1061
rect 1586 1058 1622 1061
rect 1698 1058 1718 1061
rect 1786 1058 1905 1061
rect 2026 1058 2086 1061
rect 2154 1058 2174 1061
rect 2178 1058 2182 1061
rect 2194 1058 2222 1061
rect 2270 1061 2273 1068
rect 2454 1062 2457 1068
rect 2226 1058 2273 1061
rect 2362 1058 2422 1061
rect 2490 1058 2494 1061
rect 2538 1058 2558 1061
rect 2578 1058 2582 1061
rect 2610 1058 2622 1061
rect 2642 1058 2646 1061
rect 2654 1061 2657 1068
rect 3550 1062 3553 1068
rect 3558 1062 3561 1068
rect 3614 1062 3617 1068
rect 2654 1058 2769 1061
rect 2802 1058 2806 1061
rect 2818 1058 2838 1061
rect 2890 1058 2918 1061
rect 2962 1058 3046 1061
rect 3066 1058 3070 1061
rect 3082 1058 3102 1061
rect 3202 1058 3206 1061
rect 3210 1058 3233 1061
rect 3242 1058 3286 1061
rect 3306 1058 3310 1061
rect 3378 1058 3406 1061
rect 3410 1058 3438 1061
rect 3442 1058 3526 1061
rect 3650 1058 3710 1061
rect 302 1052 305 1058
rect 1526 1052 1529 1058
rect -26 1051 -22 1052
rect -26 1048 6 1051
rect 314 1048 318 1051
rect 514 1048 678 1051
rect 906 1048 966 1051
rect 970 1048 990 1051
rect 1130 1048 1206 1051
rect 1210 1048 1214 1051
rect 1354 1048 1358 1051
rect 1378 1048 1406 1051
rect 1426 1048 1470 1051
rect 1498 1048 1526 1051
rect 1538 1048 1654 1051
rect 1666 1048 1726 1051
rect 1778 1048 1894 1051
rect 1902 1051 1905 1058
rect 1902 1048 2022 1051
rect 2030 1048 2078 1051
rect 2122 1048 2262 1051
rect 2314 1048 2369 1051
rect 2442 1048 2446 1051
rect 2566 1051 2569 1058
rect 2766 1052 2769 1058
rect 3230 1052 3233 1058
rect 3286 1052 3289 1058
rect 2506 1048 2569 1051
rect 2634 1048 2694 1051
rect 2714 1048 2726 1051
rect 2738 1048 2750 1051
rect 2794 1048 2806 1051
rect 2834 1048 2998 1051
rect 3018 1048 3094 1051
rect 3114 1048 3142 1051
rect 3354 1048 3390 1051
rect 3398 1048 3454 1051
rect 3490 1048 3494 1051
rect 3514 1048 3665 1051
rect 678 1042 681 1048
rect 2030 1042 2033 1048
rect 2102 1042 2105 1048
rect 2366 1042 2369 1048
rect 3102 1042 3105 1048
rect 458 1038 486 1041
rect 890 1038 926 1041
rect 1098 1038 1422 1041
rect 1498 1038 1510 1041
rect 1514 1038 1574 1041
rect 1634 1038 1990 1041
rect 2562 1038 2590 1041
rect 2594 1038 2758 1041
rect 2866 1038 2870 1041
rect 3398 1041 3401 1048
rect 3662 1042 3665 1048
rect 3138 1038 3401 1041
rect 3410 1038 3478 1041
rect 3482 1038 3502 1041
rect 3594 1038 3614 1041
rect 3626 1038 3646 1041
rect 442 1028 630 1031
rect 1138 1028 1150 1031
rect 1354 1028 1758 1031
rect 1770 1028 1822 1031
rect 2126 1031 2129 1038
rect 1842 1028 2129 1031
rect 2234 1028 2838 1031
rect 2934 1031 2937 1038
rect 2934 1028 3022 1031
rect 3170 1028 3214 1031
rect 3226 1028 3262 1031
rect 3266 1028 3294 1031
rect 3346 1028 3398 1031
rect 3402 1028 3510 1031
rect 3610 1028 3614 1031
rect 3630 1028 3718 1031
rect 3030 1022 3033 1028
rect 3630 1022 3633 1028
rect 266 1018 486 1021
rect 1106 1018 1646 1021
rect 1650 1018 1710 1021
rect 1722 1018 2062 1021
rect 2138 1018 2150 1021
rect 2366 1018 2918 1021
rect 2938 1018 3014 1021
rect 3042 1018 3046 1021
rect 3050 1018 3054 1021
rect 3202 1018 3486 1021
rect 3658 1018 3710 1021
rect 2366 1012 2369 1018
rect 1170 1008 1278 1011
rect 1434 1008 1630 1011
rect 1642 1008 1646 1011
rect 1714 1008 2366 1011
rect 2434 1008 2462 1011
rect 2466 1008 2750 1011
rect 2754 1008 3318 1011
rect 344 1003 346 1007
rect 350 1003 353 1007
rect 358 1003 360 1007
rect 422 1002 425 1008
rect 1360 1003 1362 1007
rect 1366 1003 1369 1007
rect 1374 1003 1376 1007
rect 2384 1003 2386 1007
rect 2390 1003 2393 1007
rect 2398 1003 2400 1007
rect 3408 1003 3410 1007
rect 3414 1003 3417 1007
rect 3422 1003 3424 1007
rect 954 998 998 1001
rect 1242 998 1254 1001
rect 1402 998 1550 1001
rect 1586 998 1590 1001
rect 1674 998 1686 1001
rect 1762 998 1854 1001
rect 1858 998 1974 1001
rect 1986 998 2158 1001
rect 2186 998 2198 1001
rect 2570 998 2726 1001
rect 2746 998 2774 1001
rect 2938 998 2950 1001
rect 2994 998 3070 1001
rect 3170 998 3174 1001
rect 3530 998 3638 1001
rect 3642 998 3694 1001
rect 242 988 390 991
rect 574 991 577 998
rect 554 988 577 991
rect 1210 988 2790 991
rect 2794 988 3294 991
rect 3314 988 3510 991
rect 3574 988 3662 991
rect 122 978 241 981
rect 306 978 390 981
rect 1266 978 1454 981
rect 1562 978 1646 981
rect 1650 978 1782 981
rect 1786 978 2118 981
rect 2162 978 2166 981
rect 2190 978 2198 981
rect 2202 978 2222 981
rect 2346 978 2470 981
rect 2494 978 2574 981
rect 2674 978 2990 981
rect 3034 978 3038 981
rect 3046 978 3054 981
rect 3058 978 3078 981
rect 3146 978 3422 981
rect 3574 981 3577 988
rect 3498 978 3577 981
rect 3586 978 3606 981
rect 238 972 241 978
rect 338 968 497 971
rect 962 968 1638 971
rect 1642 968 1782 971
rect 1858 968 1910 971
rect 1914 968 1958 971
rect 1970 968 2230 971
rect 2294 971 2297 978
rect 2494 972 2497 978
rect 2294 968 2390 971
rect 2394 968 2494 971
rect 2602 968 2782 971
rect 2890 968 2926 971
rect 2954 968 2958 971
rect 3018 968 3078 971
rect 3082 968 3086 971
rect 3162 968 3182 971
rect 3474 968 3502 971
rect 3506 968 3566 971
rect 3594 968 3646 971
rect 3650 968 3689 971
rect 326 961 329 968
rect 494 962 497 968
rect 2558 962 2561 968
rect 2566 962 2569 968
rect 3150 962 3153 968
rect 3230 962 3233 968
rect 3366 962 3369 968
rect 3686 962 3689 968
rect 298 958 329 961
rect 474 958 478 961
rect 650 958 1102 961
rect 1154 958 1198 961
rect 1602 958 1606 961
rect 1626 958 1654 961
rect 1690 958 1718 961
rect 1746 958 1766 961
rect 1770 958 1958 961
rect 1978 958 2118 961
rect 2154 958 2190 961
rect 2194 958 2270 961
rect 2274 958 2286 961
rect 2394 958 2478 961
rect 2650 958 2686 961
rect 2690 958 2718 961
rect 2722 958 2830 961
rect 2842 958 2846 961
rect 2914 958 2942 961
rect 2946 958 3150 961
rect 3154 958 3198 961
rect 3234 958 3246 961
rect 3386 958 3478 961
rect 3490 958 3497 961
rect 2342 952 2345 958
rect 322 948 334 951
rect 474 948 478 951
rect 706 948 750 951
rect 810 948 910 951
rect 1034 948 1166 951
rect 1338 948 1390 951
rect 1450 948 1550 951
rect 1570 948 1694 951
rect 1722 948 1726 951
rect 1770 948 1806 951
rect 1826 948 1830 951
rect 1890 948 1910 951
rect 1922 948 1926 951
rect 1954 948 1982 951
rect 2170 948 2174 951
rect 2210 948 2278 951
rect 2290 948 2313 951
rect 2354 948 2366 951
rect 2382 951 2385 958
rect 2526 952 2529 958
rect 2534 952 2537 958
rect 2582 952 2585 958
rect 2378 948 2385 951
rect 2418 948 2422 951
rect 2482 948 2502 951
rect 2626 948 2630 951
rect 2658 948 2662 951
rect 2690 948 2702 951
rect 2738 948 2742 951
rect 2770 948 2806 951
rect 2810 948 2814 951
rect 2842 948 2846 951
rect 2874 948 2878 951
rect 2930 948 2966 951
rect 2978 948 2982 951
rect 2994 948 2998 951
rect 3058 948 3062 951
rect 3090 948 3118 951
rect 3130 948 3134 951
rect 3146 948 3254 951
rect 3258 948 3262 951
rect 3298 948 3310 951
rect 3338 948 3358 951
rect 3362 948 3398 951
rect 3478 948 3486 951
rect 3494 951 3497 958
rect 3546 958 3550 961
rect 3626 958 3630 961
rect 3634 958 3670 961
rect 3690 958 3758 961
rect 3510 952 3513 958
rect 3494 948 3502 951
rect 3530 948 3774 951
rect 310 942 313 948
rect 670 942 673 948
rect 2054 942 2057 948
rect 2310 942 2313 948
rect 3006 942 3009 948
rect 274 938 286 941
rect 394 938 454 941
rect 490 938 534 941
rect 794 938 830 941
rect 834 938 950 941
rect 1010 938 1046 941
rect 1146 938 1182 941
rect 1186 938 1398 941
rect 1426 938 1494 941
rect 1498 938 1542 941
rect 1562 938 1566 941
rect 1594 938 1598 941
rect 1602 938 1758 941
rect 1810 938 1814 941
rect 1850 938 1854 941
rect 1866 938 1950 941
rect 2182 938 2262 941
rect 2282 938 2302 941
rect 2338 938 2438 941
rect 2490 938 2510 941
rect 2574 938 2582 941
rect 2586 938 2598 941
rect 2666 938 2678 941
rect 2746 938 2801 941
rect 2810 938 2838 941
rect 2866 938 2998 941
rect 3066 938 3070 941
rect 3178 938 3190 941
rect 3274 938 3278 941
rect 3306 938 3350 941
rect 3478 941 3481 948
rect 3526 942 3529 948
rect 3370 938 3481 941
rect 3490 938 3518 941
rect 3570 938 3726 941
rect 106 928 334 931
rect 410 928 430 931
rect 434 928 446 931
rect 514 928 537 931
rect 602 928 657 931
rect 534 922 537 928
rect 654 922 657 928
rect 1598 931 1601 938
rect 1546 928 1601 931
rect 1634 928 1662 931
rect 1666 928 1686 931
rect 1706 928 1710 931
rect 1806 931 1809 938
rect 1738 928 1809 931
rect 1838 931 1841 938
rect 1838 928 1966 931
rect 1974 931 1977 938
rect 2182 931 2185 938
rect 1974 928 2185 931
rect 2202 928 2206 931
rect 2226 928 2350 931
rect 2362 928 2390 931
rect 2478 931 2481 938
rect 2458 928 2481 931
rect 2534 932 2537 938
rect 2646 932 2649 938
rect 2686 932 2689 938
rect 2798 932 2801 938
rect 2618 928 2622 931
rect 2834 928 2854 931
rect 2866 928 2926 931
rect 2970 928 3030 931
rect 3122 928 3134 931
rect 3170 928 3182 931
rect 3186 928 3246 931
rect 3266 928 3270 931
rect 3290 928 3446 931
rect 3562 928 3622 931
rect 3722 928 3750 931
rect 1046 922 1049 928
rect 18 918 46 921
rect 410 918 422 921
rect 1458 918 1726 921
rect 1734 918 2182 921
rect 2242 918 2630 921
rect 2646 921 2649 928
rect 2646 918 2814 921
rect 2818 918 2990 921
rect 3026 918 3086 921
rect 3246 921 3249 928
rect 3510 922 3513 928
rect 3670 922 3673 928
rect 3246 918 3358 921
rect 3578 918 3590 921
rect 1734 912 1737 918
rect 130 908 238 911
rect 242 908 822 911
rect 1194 908 1222 911
rect 1226 908 1294 911
rect 1314 908 1734 911
rect 1802 908 1830 911
rect 1922 908 2062 911
rect 2074 908 2078 911
rect 2122 908 2174 911
rect 2178 908 2190 911
rect 2258 908 2294 911
rect 2322 908 2374 911
rect 2418 908 2518 911
rect 2562 908 2582 911
rect 2594 908 2710 911
rect 2874 908 2894 911
rect 2962 908 3294 911
rect 3474 908 3582 911
rect 3666 908 3686 911
rect 3698 908 3710 911
rect 848 903 850 907
rect 854 903 857 907
rect 862 903 864 907
rect 1880 903 1882 907
rect 1886 903 1889 907
rect 1894 903 1896 907
rect 2766 902 2769 908
rect 2904 903 2906 907
rect 2910 903 2913 907
rect 2918 903 2920 907
rect 122 898 174 901
rect 202 898 462 901
rect 466 898 502 901
rect 506 898 526 901
rect 1114 898 1430 901
rect 1530 898 1590 901
rect 1642 898 1830 901
rect 1850 898 1870 901
rect 1970 898 2230 901
rect 2362 898 2446 901
rect 2466 898 2486 901
rect 2538 898 2558 901
rect 2562 898 2614 901
rect 2834 898 2870 901
rect 3034 898 3102 901
rect 3162 898 3230 901
rect 3298 898 3526 901
rect 314 888 318 891
rect 402 888 406 891
rect 418 888 430 891
rect 458 888 462 891
rect 498 888 526 891
rect 530 888 537 891
rect 554 888 574 891
rect 938 888 958 891
rect 1226 888 1310 891
rect 1322 888 1598 891
rect 1602 888 1609 891
rect 1786 888 1838 891
rect 1862 888 1870 891
rect 1874 888 1894 891
rect 1906 888 1926 891
rect 1962 888 1966 891
rect 1970 888 2254 891
rect 2266 888 2310 891
rect 2410 888 2438 891
rect 2526 888 3046 891
rect 3098 888 3126 891
rect 3130 888 3166 891
rect 3522 888 3558 891
rect 86 882 89 888
rect 210 878 214 881
rect 334 881 337 888
rect 334 878 382 881
rect 386 878 446 881
rect 450 878 470 881
rect 474 878 534 881
rect 538 878 558 881
rect 590 881 593 888
rect 578 878 686 881
rect 742 881 745 888
rect 690 878 745 881
rect 1006 882 1009 888
rect 1198 881 1201 888
rect 2526 882 2529 888
rect 3302 882 3305 888
rect 3406 882 3409 888
rect 1122 878 1201 881
rect 1290 878 1294 881
rect 1314 878 1417 881
rect 1458 878 1558 881
rect 1562 878 1678 881
rect 1722 878 1742 881
rect 1770 878 1774 881
rect 1802 878 1910 881
rect 2234 878 2342 881
rect 2370 878 2374 881
rect 2426 878 2430 881
rect 2482 878 2502 881
rect 2506 878 2526 881
rect 2610 878 2638 881
rect 2690 878 2702 881
rect 2770 878 2830 881
rect 2850 878 2854 881
rect 2882 878 2886 881
rect 2890 878 2918 881
rect 2986 878 3070 881
rect 3090 878 3094 881
rect 3210 878 3294 881
rect 3322 878 3326 881
rect 3378 878 3382 881
rect 3450 878 3582 881
rect 3642 878 3654 881
rect 1022 872 1025 878
rect 1414 872 1417 878
rect 2750 872 2753 878
rect 70 868 278 871
rect 306 868 502 871
rect 506 868 646 871
rect 650 868 654 871
rect 858 868 902 871
rect 1146 868 1150 871
rect 1154 868 1206 871
rect 1274 868 1278 871
rect 1418 868 1486 871
rect 1506 868 1510 871
rect 1538 868 1590 871
rect 1666 868 1710 871
rect 1778 868 1782 871
rect 1946 868 1974 871
rect 2114 868 2174 871
rect 2182 868 2486 871
rect 2498 868 2502 871
rect 2522 868 2582 871
rect 2618 868 2622 871
rect 2634 868 2662 871
rect 2698 868 2734 871
rect 2842 868 2846 871
rect 2858 868 2870 871
rect 2906 868 2910 871
rect 2922 868 2934 871
rect 2958 871 2961 878
rect 3030 872 3033 878
rect 2954 868 2961 871
rect 2970 868 2974 871
rect 3010 868 3017 871
rect 3106 868 3142 871
rect 3162 868 3198 871
rect 3246 868 3262 871
rect 3330 868 3342 871
rect 3410 868 3454 871
rect 3514 868 3590 871
rect 3626 868 3638 871
rect 3666 868 3686 871
rect 3706 868 3718 871
rect 3722 868 3729 871
rect 70 862 73 868
rect 1094 862 1097 868
rect 1126 862 1129 868
rect 1134 862 1137 868
rect 1870 862 1873 868
rect 2054 862 2057 868
rect 330 858 342 861
rect 378 858 398 861
rect 434 858 478 861
rect 1082 858 1086 861
rect 1202 858 1230 861
rect 1274 858 1350 861
rect 1522 858 1574 861
rect 1602 858 1614 861
rect 1650 858 1670 861
rect 1698 858 1774 861
rect 1922 858 1966 861
rect 2182 861 2185 868
rect 2146 858 2185 861
rect 2418 858 2430 861
rect 2434 858 2454 861
rect 2458 858 2622 861
rect 2670 861 2673 868
rect 2650 858 2673 861
rect 2678 862 2681 868
rect 2694 862 2697 868
rect 2814 862 2817 868
rect 3014 862 3017 868
rect 3246 862 3249 868
rect 2770 858 2774 861
rect 2786 858 2790 861
rect 2818 858 2990 861
rect 3106 858 3110 861
rect 3114 858 3166 861
rect 3210 858 3214 861
rect 3338 858 3350 861
rect 3354 858 3462 861
rect 3466 858 3478 861
rect 3482 858 3566 861
rect 3570 858 3670 861
rect 3698 858 3742 861
rect 234 848 406 851
rect 1186 848 1206 851
rect 1306 848 1414 851
rect 1418 848 1513 851
rect 1510 842 1513 848
rect 1526 848 1566 851
rect 1570 848 1574 851
rect 1626 848 1630 851
rect 1634 848 1718 851
rect 1730 848 1750 851
rect 1754 848 1790 851
rect 1810 848 1814 851
rect 1834 848 1878 851
rect 1938 848 1998 851
rect 2034 848 2038 851
rect 2382 848 2406 851
rect 2434 848 2462 851
rect 2658 848 2937 851
rect 2962 848 3070 851
rect 3118 848 3161 851
rect 1526 842 1529 848
rect 2382 842 2385 848
rect 2934 842 2937 848
rect 3118 842 3121 848
rect 3158 842 3161 848
rect 3210 848 3254 851
rect 3346 848 3358 851
rect 3386 848 3449 851
rect 3458 848 3470 851
rect 3482 848 3518 851
rect 3562 848 3574 851
rect 3634 848 3638 851
rect 186 838 262 841
rect 378 838 422 841
rect 1154 838 1470 841
rect 1618 838 1814 841
rect 1818 838 1902 841
rect 1954 838 1982 841
rect 1986 838 2126 841
rect 2514 838 2542 841
rect 2546 838 2702 841
rect 2770 838 2806 841
rect 2858 838 2894 841
rect 2898 838 2902 841
rect 2970 838 2982 841
rect 2986 838 3006 841
rect 3058 838 3070 841
rect 3174 841 3177 848
rect 3446 842 3449 848
rect 3174 838 3214 841
rect 3242 838 3262 841
rect 3322 838 3350 841
rect 3354 838 3398 841
rect 3450 838 3486 841
rect 3490 838 3590 841
rect 3594 838 3702 841
rect 1942 832 1945 838
rect 42 828 958 831
rect 962 828 1398 831
rect 1434 828 1665 831
rect 1682 828 1782 831
rect 1786 828 1934 831
rect 1954 828 2361 831
rect 2370 828 2422 831
rect 2498 828 2534 831
rect 2538 828 2654 831
rect 2658 828 3070 831
rect 3086 831 3089 838
rect 3086 828 3142 831
rect 3398 831 3401 838
rect 3398 828 3598 831
rect 3602 828 3609 831
rect 3626 828 3646 831
rect 3690 828 3702 831
rect 3714 828 3734 831
rect 1662 822 1665 828
rect 170 818 174 821
rect 258 818 366 821
rect 370 818 390 821
rect 666 818 670 821
rect 738 818 910 821
rect 914 818 1294 821
rect 1298 818 1310 821
rect 1330 818 1614 821
rect 1898 818 2062 821
rect 2066 818 2118 821
rect 2138 818 2326 821
rect 2358 821 2361 828
rect 2358 818 2662 821
rect 2666 818 2758 821
rect 2802 818 3038 821
rect 3042 818 3102 821
rect 3146 818 3182 821
rect 3490 818 3518 821
rect 2134 812 2137 818
rect 498 808 510 811
rect 762 808 790 811
rect 1474 808 1630 811
rect 1634 808 1750 811
rect 1818 808 1934 811
rect 2210 808 2222 811
rect 2458 808 2462 811
rect 2490 808 2566 811
rect 2618 808 2694 811
rect 2954 808 3046 811
rect 3050 808 3150 811
rect 3154 808 3182 811
rect 3458 808 3638 811
rect 344 803 346 807
rect 350 803 353 807
rect 358 803 360 807
rect 1360 803 1362 807
rect 1366 803 1369 807
rect 1374 803 1376 807
rect 2384 803 2386 807
rect 2390 803 2393 807
rect 2398 803 2400 807
rect 3408 803 3410 807
rect 3414 803 3417 807
rect 3422 803 3424 807
rect 1170 798 1326 801
rect 1498 798 1710 801
rect 1722 798 1846 801
rect 1858 798 1862 801
rect 1874 798 2142 801
rect 2154 798 2182 801
rect 2186 798 2238 801
rect 2330 798 2374 801
rect 2498 798 2550 801
rect 2706 798 2774 801
rect 2890 798 3222 801
rect 3610 798 3686 801
rect 1258 788 2838 791
rect 2850 788 2934 791
rect 2986 788 3006 791
rect 3430 788 3438 791
rect 3442 788 3622 791
rect 3650 788 3662 791
rect 3690 788 3726 791
rect 3230 782 3233 788
rect 186 778 206 781
rect 274 778 302 781
rect 810 778 862 781
rect 1162 778 1166 781
rect 1426 778 1689 781
rect 1866 778 2150 781
rect 2178 778 2182 781
rect 2218 778 2222 781
rect 2282 778 2286 781
rect 2346 778 2358 781
rect 2362 778 2457 781
rect 2466 778 2526 781
rect 2954 778 2974 781
rect 3018 778 3094 781
rect 3370 778 3505 781
rect 3546 778 3590 781
rect 3594 778 3630 781
rect 3658 778 3670 781
rect 1686 772 1689 778
rect 2454 772 2457 778
rect 2702 772 2705 778
rect 130 768 158 771
rect 162 768 198 771
rect 202 768 310 771
rect 366 768 374 771
rect 378 768 398 771
rect 426 768 566 771
rect 802 768 838 771
rect 842 768 886 771
rect 1130 768 1254 771
rect 1458 768 1510 771
rect 1738 768 1886 771
rect 1914 768 2078 771
rect 2082 768 2294 771
rect 2306 768 2334 771
rect 2338 768 2422 771
rect 2426 768 2430 771
rect 2458 768 2526 771
rect 2530 768 2582 771
rect 2770 768 2798 771
rect 2842 768 2854 771
rect 2862 771 2865 778
rect 2862 768 2910 771
rect 2962 768 2966 771
rect 3018 768 3022 771
rect 3034 768 3054 771
rect 3094 771 3097 778
rect 3502 772 3505 778
rect 3094 768 3142 771
rect 3186 768 3230 771
rect 3506 768 3590 771
rect 3594 768 3686 771
rect 3726 771 3729 778
rect 3726 768 3750 771
rect 54 761 57 768
rect 54 758 310 761
rect 314 758 678 761
rect 826 758 838 761
rect 1034 758 1182 761
rect 1314 758 1318 761
rect 1546 758 1550 761
rect 1578 758 1582 761
rect 1602 758 1766 761
rect 1802 758 1806 761
rect 1810 758 1830 761
rect 1834 758 2262 761
rect 2266 758 2582 761
rect 2626 758 2769 761
rect 2834 758 2886 761
rect 2974 761 2977 768
rect 2906 758 2977 761
rect 3078 761 3081 768
rect 3078 758 3110 761
rect 3114 758 3134 761
rect 3178 758 3254 761
rect 3258 758 3262 761
rect 3386 758 3446 761
rect 3462 761 3465 768
rect 3462 758 3486 761
rect 3546 758 3550 761
rect 3610 758 3766 761
rect 3770 758 3774 761
rect 1510 752 1513 758
rect 74 748 78 751
rect 138 748 166 751
rect 242 748 270 751
rect 290 748 294 751
rect 306 748 486 751
rect 786 748 790 751
rect 834 748 886 751
rect 1122 748 1174 751
rect 1194 748 1222 751
rect 1522 748 1550 751
rect 1570 748 1574 751
rect 1642 748 1678 751
rect 1754 748 1758 751
rect 2058 748 2094 751
rect 2130 748 2230 751
rect 2266 748 2326 751
rect 2330 748 2430 751
rect 2486 748 2494 751
rect 2514 748 2518 751
rect 2570 748 2686 751
rect 2698 748 2702 751
rect 2730 748 2758 751
rect 2766 751 2769 758
rect 2766 748 2833 751
rect 106 738 150 741
rect 214 741 217 748
rect 454 742 457 748
rect 214 738 230 741
rect 466 738 486 741
rect 490 738 502 741
rect 774 741 777 748
rect 562 738 641 741
rect 774 738 822 741
rect 826 738 902 741
rect 1170 738 1230 741
rect 1514 738 1542 741
rect 1674 738 1806 741
rect 1810 738 1814 741
rect 1818 738 1950 741
rect 1990 741 1993 748
rect 2830 742 2833 748
rect 2882 748 2918 751
rect 2922 748 2926 751
rect 2994 748 3014 751
rect 3058 748 3278 751
rect 3338 748 3361 751
rect 3394 748 3478 751
rect 3582 751 3585 758
rect 3514 748 3598 751
rect 3658 748 3670 751
rect 3690 748 3758 751
rect 2854 742 2857 748
rect 3358 742 3361 748
rect 1990 738 2086 741
rect 2122 738 2158 741
rect 2178 738 2286 741
rect 2290 738 2406 741
rect 2426 738 2478 741
rect 2490 738 2494 741
rect 2626 738 2734 741
rect 2754 738 2798 741
rect 2938 738 2958 741
rect 2962 738 2982 741
rect 3002 738 3022 741
rect 3090 738 3190 741
rect 3194 738 3206 741
rect 3250 738 3262 741
rect 3306 738 3310 741
rect 3402 738 3470 741
rect 3578 738 3710 741
rect 638 732 641 738
rect 82 728 150 731
rect 154 728 246 731
rect 250 728 278 731
rect 322 728 342 731
rect 346 728 390 731
rect 394 728 470 731
rect 658 728 734 731
rect 738 728 1006 731
rect 1046 731 1049 738
rect 1046 728 1150 731
rect 1270 731 1273 738
rect 1226 728 1273 731
rect 1610 728 1630 731
rect 1714 728 1742 731
rect 1974 731 1977 738
rect 2454 732 2457 738
rect 1754 728 1977 731
rect 2002 728 2078 731
rect 2082 728 2198 731
rect 2378 728 2382 731
rect 2410 728 2438 731
rect 2474 728 2478 731
rect 2490 728 2630 731
rect 2674 728 2678 731
rect 2690 728 2726 731
rect 2778 728 2814 731
rect 2862 731 2865 738
rect 2818 728 2865 731
rect 2898 728 2934 731
rect 2954 728 2966 731
rect 2986 728 3014 731
rect 3054 731 3057 738
rect 3050 728 3057 731
rect 3062 732 3065 738
rect 3114 728 3118 731
rect 3122 728 3206 731
rect 3234 728 3246 731
rect 3298 728 3305 731
rect 622 722 625 728
rect 106 718 214 721
rect 218 718 225 721
rect 250 718 262 721
rect 270 718 422 721
rect 754 718 1150 721
rect 1502 721 1505 728
rect 3302 722 3305 728
rect 3378 728 3422 731
rect 3450 728 3454 731
rect 3502 731 3505 738
rect 3502 728 3614 731
rect 3626 728 3686 731
rect 3318 722 3321 728
rect 3334 722 3337 728
rect 3462 722 3465 728
rect 3710 722 3713 728
rect 1466 718 1505 721
rect 1514 718 1758 721
rect 1778 718 3073 721
rect 3082 718 3126 721
rect 3138 718 3158 721
rect 3162 718 3169 721
rect 3178 718 3182 721
rect 3378 718 3382 721
rect 3558 718 3574 721
rect 3650 718 3670 721
rect 270 711 273 718
rect 234 708 273 711
rect 410 708 462 711
rect 594 708 606 711
rect 610 708 702 711
rect 794 708 830 711
rect 1122 708 1238 711
rect 1298 708 1358 711
rect 1362 708 1542 711
rect 1922 708 2222 711
rect 2226 708 2406 711
rect 2410 708 2814 711
rect 2842 708 2862 711
rect 2930 708 3038 711
rect 3070 711 3073 718
rect 3070 708 3254 711
rect 3558 711 3561 718
rect 3614 712 3617 718
rect 3322 708 3561 711
rect 3570 708 3598 711
rect 3602 708 3606 711
rect 3682 708 3718 711
rect 848 703 850 707
rect 854 703 857 707
rect 862 703 864 707
rect 1880 703 1882 707
rect 1886 703 1889 707
rect 1894 703 1896 707
rect 2904 703 2906 707
rect 2910 703 2913 707
rect 2918 703 2920 707
rect 74 698 86 701
rect 170 698 254 701
rect 410 698 582 701
rect 666 698 838 701
rect 962 698 1502 701
rect 1538 698 1670 701
rect 1690 698 1718 701
rect 2162 698 2174 701
rect 2202 698 2302 701
rect 2450 698 2510 701
rect 2666 698 2726 701
rect 2730 698 2750 701
rect 2826 698 2846 701
rect 2858 698 2894 701
rect 2994 698 3214 701
rect 3298 698 3510 701
rect 3514 698 3558 701
rect 3578 698 3622 701
rect 3634 698 3758 701
rect 314 688 326 691
rect 330 688 382 691
rect 978 688 1046 691
rect 1402 688 1478 691
rect 1482 688 1494 691
rect 1570 688 1598 691
rect 1890 688 1966 691
rect 2066 688 2118 691
rect 2258 688 2278 691
rect 2322 688 2438 691
rect 2450 688 2470 691
rect 2482 688 2534 691
rect 2738 688 2774 691
rect 2810 688 2854 691
rect 2870 688 2878 691
rect 2882 688 2894 691
rect 2902 688 2910 691
rect 2914 688 2998 691
rect 3082 688 3110 691
rect 3298 688 3310 691
rect 3350 688 3478 691
rect 3490 688 3542 691
rect 3626 688 3750 691
rect 86 682 89 688
rect 178 678 190 681
rect 194 678 198 681
rect 238 681 241 688
rect 238 678 326 681
rect 330 678 358 681
rect 422 681 425 688
rect 418 678 425 681
rect 450 678 489 681
rect 498 678 718 681
rect 974 681 977 688
rect 1150 682 1153 688
rect 1742 682 1745 688
rect 722 678 977 681
rect 1282 678 1318 681
rect 1346 678 1374 681
rect 1410 678 1462 681
rect 1578 678 1622 681
rect 1946 678 1966 681
rect 1970 678 1974 681
rect 1986 678 2046 681
rect 2174 681 2177 688
rect 2294 682 2297 688
rect 2050 678 2262 681
rect 2354 678 2366 681
rect 2450 678 2470 681
rect 2474 678 2502 681
rect 2642 678 2686 681
rect 2762 678 2838 681
rect 2874 678 2926 681
rect 2930 678 2998 681
rect 3010 678 3158 681
rect 3262 681 3265 688
rect 3218 678 3286 681
rect 3350 681 3353 688
rect 3290 678 3353 681
rect 3362 678 3366 681
rect 3402 678 3422 681
rect 3506 678 3510 681
rect 3606 681 3609 688
rect 3514 678 3609 681
rect 3714 678 3758 681
rect 486 672 489 678
rect 210 668 238 671
rect 282 668 374 671
rect 378 668 398 671
rect 418 668 422 671
rect 458 668 470 671
rect 530 668 534 671
rect 1134 671 1137 678
rect 1262 671 1265 678
rect 1494 672 1497 678
rect 1134 668 1265 671
rect 1314 668 1342 671
rect 1418 668 1422 671
rect 1522 668 1566 671
rect 1602 668 1606 671
rect 1726 671 1729 678
rect 1726 668 1862 671
rect 1962 668 2022 671
rect 2058 668 2254 671
rect 2282 668 2286 671
rect 2290 668 2417 671
rect 2474 668 2486 671
rect 2530 668 2710 671
rect 2778 668 2782 671
rect 2786 668 2886 671
rect 2890 668 3094 671
rect 3098 668 3102 671
rect 3282 668 3534 671
rect 3538 668 3598 671
rect 3602 668 3726 671
rect 582 662 585 668
rect 638 662 641 668
rect 1926 662 1929 668
rect 1950 662 1953 668
rect 210 658 214 661
rect 394 658 398 661
rect 402 658 422 661
rect 482 658 526 661
rect 1018 658 1078 661
rect 1242 658 1246 661
rect 1250 658 1286 661
rect 1410 658 1438 661
rect 1442 658 1614 661
rect 1618 658 1654 661
rect 1970 658 1990 661
rect 2034 658 2038 661
rect 2098 658 2102 661
rect 2130 658 2142 661
rect 2178 658 2182 661
rect 2234 658 2246 661
rect 2250 658 2262 661
rect 2338 658 2342 661
rect 2362 658 2406 661
rect 2414 661 2417 668
rect 3118 662 3121 668
rect 2414 658 2662 661
rect 2666 658 2742 661
rect 2746 658 2790 661
rect 2794 658 2846 661
rect 2850 658 2974 661
rect 3002 658 3006 661
rect 3042 658 3046 661
rect 3162 658 3166 661
rect 3202 658 3206 661
rect 3242 658 3310 661
rect 3338 658 3374 661
rect 3378 658 3398 661
rect 3442 658 3558 661
rect 3570 658 3590 661
rect 3666 658 3670 661
rect 3686 658 3742 661
rect 3686 652 3689 658
rect 402 648 558 651
rect 898 648 974 651
rect 1242 648 1310 651
rect 1330 648 1350 651
rect 1354 648 1454 651
rect 1514 648 1638 651
rect 1666 648 1726 651
rect 1850 648 1886 651
rect 1938 648 1974 651
rect 1978 648 1990 651
rect 1994 648 1998 651
rect 2010 648 2014 651
rect 2194 648 2302 651
rect 2314 648 2350 651
rect 2370 648 2470 651
rect 2498 648 2502 651
rect 2586 648 3174 651
rect 3178 648 3222 651
rect 3286 648 3326 651
rect 3482 648 3518 651
rect 3562 648 3574 651
rect 3586 648 3686 651
rect 3730 648 3750 651
rect 3762 648 3766 651
rect 3286 642 3289 648
rect 1266 638 1366 641
rect 1634 638 1694 641
rect 1698 638 1854 641
rect 1858 638 1910 641
rect 1954 638 2054 641
rect 2138 638 2246 641
rect 2250 638 2318 641
rect 2490 638 2510 641
rect 2514 638 2758 641
rect 2762 638 2774 641
rect 2786 638 2790 641
rect 2802 638 2830 641
rect 2882 638 2886 641
rect 2906 638 2910 641
rect 2978 638 2990 641
rect 3018 638 3062 641
rect 3146 638 3254 641
rect 3258 638 3270 641
rect 3706 638 3750 641
rect 3678 632 3681 638
rect 1282 628 1334 631
rect 1338 628 1614 631
rect 1618 628 1710 631
rect 1890 628 1942 631
rect 1946 628 2006 631
rect 2258 628 3102 631
rect 3114 628 3342 631
rect 3386 628 3454 631
rect 3458 628 3638 631
rect 722 618 889 621
rect 1066 618 1590 621
rect 1834 618 1838 621
rect 1842 618 2166 621
rect 2170 618 2254 621
rect 2278 618 2286 621
rect 2290 618 2366 621
rect 2378 618 3462 621
rect 3466 618 3510 621
rect 3602 618 3694 621
rect 874 608 878 611
rect 886 611 889 618
rect 886 608 1174 611
rect 1258 608 1286 611
rect 1578 608 2014 611
rect 2026 608 2086 611
rect 2138 608 2198 611
rect 2210 608 2214 611
rect 2274 608 2318 611
rect 2498 608 2622 611
rect 2726 608 2766 611
rect 2778 608 2942 611
rect 3162 608 3190 611
rect 3314 608 3390 611
rect 3434 608 3454 611
rect 3458 608 3510 611
rect 3658 608 3686 611
rect 344 603 346 607
rect 350 603 353 607
rect 358 603 360 607
rect 1360 603 1362 607
rect 1366 603 1369 607
rect 1374 603 1376 607
rect 2384 603 2386 607
rect 2390 603 2393 607
rect 2398 603 2400 607
rect 2726 602 2729 608
rect 3408 603 3410 607
rect 3414 603 3417 607
rect 3422 603 3424 607
rect 818 598 1238 601
rect 1442 598 1454 601
rect 1506 598 1622 601
rect 1626 598 1654 601
rect 1698 598 2086 601
rect 2098 598 2142 601
rect 2146 598 2238 601
rect 2442 598 2486 601
rect 2538 598 2582 601
rect 2586 598 2713 601
rect 2722 598 2726 601
rect 2746 598 2878 601
rect 2882 598 3118 601
rect 3186 598 3286 601
rect 3290 598 3342 601
rect 3674 598 3702 601
rect 282 588 310 591
rect 514 588 542 591
rect 842 588 1382 591
rect 1394 588 1486 591
rect 1594 588 1598 591
rect 1754 588 1782 591
rect 2066 588 2070 591
rect 2326 591 2329 598
rect 2090 588 2366 591
rect 2378 588 2446 591
rect 2522 588 2526 591
rect 2710 591 2713 598
rect 2710 588 2726 591
rect 2730 588 3454 591
rect 210 578 230 581
rect 554 578 974 581
rect 1146 578 1486 581
rect 1490 578 1534 581
rect 1722 578 3110 581
rect 3122 578 3177 581
rect 3258 578 3382 581
rect 3674 578 3734 581
rect 3174 572 3177 578
rect 370 568 398 571
rect 402 568 438 571
rect 450 568 510 571
rect 562 568 630 571
rect 1058 568 1142 571
rect 1146 568 1150 571
rect 1162 568 1246 571
rect 1306 568 1310 571
rect 1314 568 1406 571
rect 1610 568 2262 571
rect 2266 568 2766 571
rect 2802 568 2822 571
rect 2890 568 2926 571
rect 2938 568 2958 571
rect 3002 568 3118 571
rect 3242 568 3334 571
rect 3570 568 3598 571
rect 3602 568 3766 571
rect 214 561 217 568
rect 214 558 238 561
rect 246 561 249 568
rect 366 562 369 568
rect 782 562 785 568
rect 3214 562 3217 568
rect 246 558 286 561
rect 426 558 502 561
rect 1138 558 1206 561
rect 1210 558 1350 561
rect 1394 558 1430 561
rect 1642 558 1646 561
rect 1842 558 2014 561
rect 2026 558 2110 561
rect 2114 558 2158 561
rect 2170 558 2230 561
rect 2242 558 2254 561
rect 2258 558 2302 561
rect 2338 558 2446 561
rect 2690 558 2694 561
rect 2710 558 2718 561
rect 2722 558 2761 561
rect 2770 558 2846 561
rect 2858 558 2870 561
rect 2962 558 2966 561
rect 2994 558 3014 561
rect 3034 558 3054 561
rect 3098 558 3142 561
rect 3186 558 3190 561
rect 3258 558 3302 561
rect 3602 558 3614 561
rect 3618 558 3646 561
rect 3650 558 3678 561
rect 282 548 462 551
rect 466 548 518 551
rect 594 548 734 551
rect 770 548 846 551
rect 1010 548 1126 551
rect 1130 548 1142 551
rect 1186 548 1214 551
rect 1298 548 1313 551
rect 1322 548 1326 551
rect 1370 548 1390 551
rect 1442 548 1566 551
rect 1602 548 1614 551
rect 1626 548 1694 551
rect 1698 548 1886 551
rect 2050 548 2246 551
rect 2250 548 2462 551
rect 2466 548 2510 551
rect 2514 548 2590 551
rect 2706 548 2710 551
rect 2722 548 2742 551
rect 2758 551 2761 558
rect 3158 552 3161 558
rect 2758 548 2774 551
rect 2874 548 2886 551
rect 2922 548 2934 551
rect 2946 548 2974 551
rect 3018 548 3126 551
rect 3170 548 3174 551
rect 3178 548 3206 551
rect 3214 548 3350 551
rect 3434 548 3438 551
rect 3470 551 3473 558
rect 3442 548 3473 551
rect 3498 548 3502 551
rect 3522 548 3534 551
rect 3554 548 3558 551
rect 3578 548 3606 551
rect 3698 548 3710 551
rect 182 541 185 548
rect 902 542 905 548
rect 1310 542 1313 548
rect 2622 542 2625 548
rect 3214 542 3217 548
rect 182 538 230 541
rect 274 538 278 541
rect 370 538 390 541
rect 434 538 486 541
rect 518 538 526 541
rect 530 538 649 541
rect 1074 538 1110 541
rect 1114 538 1118 541
rect 1226 538 1262 541
rect 1314 538 1366 541
rect 1418 538 1446 541
rect 1466 538 1470 541
rect 1514 538 1542 541
rect 646 532 649 538
rect 1030 532 1033 538
rect 1550 532 1553 541
rect 1562 538 1638 541
rect 1690 538 1710 541
rect 1806 538 1918 541
rect 1954 538 2078 541
rect 2082 538 2134 541
rect 2210 538 2278 541
rect 2522 538 2526 541
rect 2698 538 2734 541
rect 2746 538 2798 541
rect 2810 538 2814 541
rect 2818 538 2998 541
rect 3074 538 3078 541
rect 3142 538 3193 541
rect 3226 538 3278 541
rect 3330 538 3342 541
rect 3514 538 3518 541
rect 3562 538 3582 541
rect 3602 538 3646 541
rect 3722 538 3745 541
rect 1806 532 1809 538
rect 2350 532 2353 538
rect 18 528 382 531
rect 410 528 414 531
rect 418 528 433 531
rect 1042 528 1078 531
rect 1114 528 1158 531
rect 1170 528 1198 531
rect 1234 528 1246 531
rect 1250 528 1390 531
rect 1442 528 1454 531
rect 1470 528 1478 531
rect 1482 528 1502 531
rect 1618 528 1622 531
rect 1650 528 1750 531
rect 1946 528 2062 531
rect 2082 528 2118 531
rect 2170 528 2214 531
rect 2354 528 2454 531
rect 2754 528 2822 531
rect 2842 528 2870 531
rect 2922 528 2926 531
rect 3086 531 3089 538
rect 3066 528 3089 531
rect 3142 532 3145 538
rect 3190 532 3193 538
rect 3274 528 3278 531
rect 3418 528 3422 531
rect 3462 531 3465 538
rect 3742 532 3745 538
rect 3450 528 3465 531
rect 3482 528 3486 531
rect 3514 528 3542 531
rect 3714 528 3721 531
rect 86 522 89 528
rect 430 522 433 528
rect 1790 522 1793 528
rect 3718 522 3721 528
rect 66 518 70 521
rect 226 518 334 521
rect 338 518 422 521
rect 634 518 918 521
rect 978 518 1102 521
rect 1170 518 1569 521
rect 1578 518 1582 521
rect 1594 518 1606 521
rect 1870 518 1982 521
rect 1986 518 2134 521
rect 2146 518 2294 521
rect 2562 518 2606 521
rect 2626 518 2774 521
rect 2810 518 2822 521
rect 2898 518 3078 521
rect 3266 518 3294 521
rect 3362 518 3406 521
rect 3538 518 3574 521
rect 3578 518 3710 521
rect 146 508 214 511
rect 258 508 422 511
rect 1018 508 1278 511
rect 1282 508 1438 511
rect 1450 508 1558 511
rect 1566 511 1569 518
rect 1566 508 1686 511
rect 1870 511 1873 518
rect 1754 508 1873 511
rect 2218 508 2894 511
rect 3026 508 3286 511
rect 3294 511 3297 518
rect 3294 508 3494 511
rect 3514 508 3630 511
rect 3634 508 3694 511
rect 3706 508 3718 511
rect 848 503 850 507
rect 854 503 857 507
rect 862 503 864 507
rect 1880 503 1882 507
rect 1886 503 1889 507
rect 1894 503 1896 507
rect 2054 502 2057 508
rect 2904 503 2906 507
rect 2910 503 2913 507
rect 2918 503 2920 507
rect 74 498 206 501
rect 370 498 382 501
rect 386 498 398 501
rect 914 498 1022 501
rect 1154 498 1270 501
rect 1354 498 1382 501
rect 1402 498 1438 501
rect 1450 498 1518 501
rect 1522 498 1686 501
rect 1690 498 1718 501
rect 1730 498 1782 501
rect 2282 498 2390 501
rect 2394 498 2446 501
rect 2458 498 2790 501
rect 2818 498 2830 501
rect 2834 498 2862 501
rect 2930 498 3038 501
rect 3042 498 3070 501
rect 3074 498 3230 501
rect 3234 498 3270 501
rect 3354 498 3398 501
rect 3658 498 3670 501
rect 3722 498 3742 501
rect 74 488 105 491
rect 178 488 222 491
rect 234 488 302 491
rect 306 488 494 491
rect 802 488 998 491
rect 1002 488 1014 491
rect 1394 488 1462 491
rect 1490 488 1590 491
rect 1726 488 1734 491
rect 1738 488 1758 491
rect 1762 488 1854 491
rect 1866 488 1918 491
rect 1922 488 1974 491
rect 2074 488 2094 491
rect 2330 488 2454 491
rect 2478 488 2790 491
rect 2818 488 2822 491
rect 2850 488 2862 491
rect 2926 491 2929 498
rect 2866 488 2929 491
rect 3106 488 3134 491
rect 3138 488 3342 491
rect 3386 488 3534 491
rect 3538 488 3542 491
rect 3706 488 3734 491
rect 102 481 105 488
rect 102 478 246 481
rect 450 478 470 481
rect 670 481 673 488
rect 1606 482 1609 488
rect 670 478 758 481
rect 762 478 806 481
rect 826 478 886 481
rect 1098 478 1126 481
rect 1346 478 1534 481
rect 1538 478 1590 481
rect 1674 478 1782 481
rect 1786 478 1798 481
rect 2170 478 2206 481
rect 2210 478 2214 481
rect 2322 478 2334 481
rect 2370 478 2382 481
rect 2418 478 2446 481
rect 2454 481 2457 488
rect 2450 478 2457 481
rect 2470 482 2473 488
rect 2478 482 2481 488
rect 2490 478 2494 481
rect 2642 478 2654 481
rect 2666 478 2718 481
rect 2722 478 2838 481
rect 2842 478 2870 481
rect 2946 478 3046 481
rect 3226 478 3238 481
rect 3306 478 3326 481
rect 3458 478 3534 481
rect 3582 481 3585 488
rect 3562 478 3585 481
rect 3670 481 3673 488
rect 3658 478 3673 481
rect 86 472 89 478
rect 178 468 286 471
rect 294 471 297 478
rect 294 468 326 471
rect 402 468 414 471
rect 422 468 462 471
rect 498 468 510 471
rect 686 468 822 471
rect 842 468 854 471
rect 858 468 870 471
rect 982 471 985 478
rect 1134 471 1137 478
rect 982 468 1137 471
rect 1142 471 1145 478
rect 1814 472 1817 478
rect 1846 472 1849 478
rect 1950 472 1953 478
rect 1142 468 1174 471
rect 1394 468 1422 471
rect 1426 468 1750 471
rect 1826 468 1833 471
rect 1898 468 1934 471
rect 2086 471 2089 478
rect 1986 468 2089 471
rect 2114 468 2142 471
rect 2158 471 2161 478
rect 2590 472 2593 478
rect 2146 468 2161 471
rect 2186 468 2494 471
rect 2498 468 2558 471
rect 2650 468 2654 471
rect 2714 468 2742 471
rect 2746 468 2769 471
rect 2778 468 2846 471
rect 2850 468 2854 471
rect 2858 468 2910 471
rect 2914 468 2974 471
rect 3194 468 3262 471
rect 3266 468 3366 471
rect 3446 471 3449 478
rect 3378 468 3449 471
rect 3462 472 3465 478
rect 3602 468 3614 471
rect 3650 468 3686 471
rect 3714 468 3734 471
rect 226 458 230 461
rect 266 458 297 461
rect 422 461 425 468
rect 686 462 689 468
rect 346 458 425 461
rect 506 458 542 461
rect 902 461 905 468
rect 818 458 905 461
rect 1082 458 1174 461
rect 1234 458 1246 461
rect 1282 458 1286 461
rect 1322 458 1382 461
rect 1422 458 1430 461
rect 1442 458 1446 461
rect 1562 458 1590 461
rect 1818 458 1838 461
rect 1858 458 1886 461
rect 1946 458 2126 461
rect 2186 458 2222 461
rect 2250 458 2254 461
rect 2266 458 2278 461
rect 2282 458 2310 461
rect 2322 458 2342 461
rect 2346 458 2358 461
rect 2362 458 2374 461
rect 2386 458 2430 461
rect 2450 458 2454 461
rect 2490 458 2502 461
rect 2506 458 2630 461
rect 2634 458 2718 461
rect 2746 458 2750 461
rect 2766 461 2769 468
rect 2766 458 2870 461
rect 2930 458 2934 461
rect 2954 458 2958 461
rect 2978 458 2982 461
rect 3026 458 3094 461
rect 3234 458 3270 461
rect 3434 458 3574 461
rect 3578 458 3590 461
rect 3594 458 3694 461
rect 3706 458 3726 461
rect 294 452 297 458
rect 242 448 262 451
rect 338 448 438 451
rect 454 451 457 458
rect 454 448 518 451
rect 826 448 838 451
rect 842 448 918 451
rect 930 448 950 451
rect 954 448 1286 451
rect 1514 448 1518 451
rect 1522 448 1526 451
rect 1562 448 1598 451
rect 1602 448 1718 451
rect 1782 451 1785 458
rect 1782 448 1910 451
rect 1914 448 1974 451
rect 2018 448 2550 451
rect 2554 448 2758 451
rect 2802 448 2838 451
rect 2850 448 2854 451
rect 2874 448 2942 451
rect 2966 448 2990 451
rect 3042 448 3046 451
rect 3218 448 3286 451
rect 3306 448 3390 451
rect 3578 448 3622 451
rect 3626 448 3654 451
rect 3658 448 3670 451
rect 266 438 318 441
rect 322 438 382 441
rect 386 438 398 441
rect 526 441 529 448
rect 514 438 529 441
rect 602 438 862 441
rect 866 438 1158 441
rect 1170 438 1190 441
rect 1194 438 1230 441
rect 1342 441 1345 448
rect 1274 438 1345 441
rect 1414 441 1417 448
rect 2966 442 2969 448
rect 1414 438 1470 441
rect 1490 438 1534 441
rect 1546 438 1886 441
rect 2090 438 2270 441
rect 2274 438 2366 441
rect 2378 438 2382 441
rect 2490 438 2494 441
rect 2538 438 2574 441
rect 2578 438 2590 441
rect 2626 438 2630 441
rect 2690 438 2694 441
rect 2826 438 2894 441
rect 3274 438 3350 441
rect 3354 438 3446 441
rect 3522 438 3582 441
rect 3618 438 3638 441
rect 558 432 561 438
rect 2646 432 2649 438
rect 1098 428 1214 431
rect 1218 428 1246 431
rect 1450 428 1734 431
rect 1746 428 1846 431
rect 1850 428 1894 431
rect 1898 428 2030 431
rect 2218 428 2230 431
rect 2442 428 2502 431
rect 2578 428 2614 431
rect 2794 428 3014 431
rect 3018 428 3022 431
rect 3138 428 3606 431
rect 3634 428 3718 431
rect 1254 421 1257 428
rect 906 418 1257 421
rect 1266 418 1478 421
rect 1602 418 1670 421
rect 2310 421 2313 428
rect 2242 418 2313 421
rect 2346 418 2526 421
rect 2530 418 2814 421
rect 2818 418 3174 421
rect 3386 418 3510 421
rect 3514 418 3558 421
rect 626 408 638 411
rect 826 408 1326 411
rect 1410 408 1502 411
rect 1610 408 1814 411
rect 1938 408 2374 411
rect 2586 408 2854 411
rect 2882 408 3254 411
rect 3258 408 3334 411
rect 3538 408 3606 411
rect 344 403 346 407
rect 350 403 353 407
rect 358 403 360 407
rect 1360 403 1362 407
rect 1366 403 1369 407
rect 1374 403 1376 407
rect 2384 403 2386 407
rect 2390 403 2393 407
rect 2398 403 2400 407
rect 3408 403 3410 407
rect 3414 403 3417 407
rect 3422 403 3424 407
rect 578 398 654 401
rect 1114 398 1350 401
rect 1466 398 1582 401
rect 1626 398 1702 401
rect 1794 398 1822 401
rect 1954 398 1990 401
rect 2130 398 2342 401
rect 2426 398 2542 401
rect 2562 398 2590 401
rect 2610 398 2742 401
rect 2794 398 2894 401
rect 2898 398 2966 401
rect 3026 398 3222 401
rect 562 388 582 391
rect 730 388 750 391
rect 922 388 1014 391
rect 1074 388 1078 391
rect 1090 388 1110 391
rect 1302 388 1478 391
rect 1582 391 1585 398
rect 1582 388 1902 391
rect 1906 388 1998 391
rect 2002 388 2134 391
rect 2194 388 2398 391
rect 2402 388 2414 391
rect 2434 388 2446 391
rect 2466 388 2582 391
rect 2634 388 2742 391
rect 2786 388 2974 391
rect 3018 388 3038 391
rect 3082 388 3102 391
rect 1302 382 1305 388
rect 978 378 1190 381
rect 1354 378 1446 381
rect 1642 378 1654 381
rect 2034 378 2038 381
rect 2050 378 2094 381
rect 2098 378 2102 381
rect 2146 378 2238 381
rect 2250 378 2366 381
rect 2378 378 2526 381
rect 2746 378 2982 381
rect 2994 378 3302 381
rect 866 368 926 371
rect 966 371 969 378
rect 946 368 1022 371
rect 1026 368 1094 371
rect 1114 368 1150 371
rect 1250 368 1742 371
rect 1870 371 1873 378
rect 1858 368 1873 371
rect 1898 368 1934 371
rect 1946 368 2033 371
rect 2098 368 2198 371
rect 2202 368 2246 371
rect 2250 368 2505 371
rect 2514 368 2518 371
rect 2522 368 2694 371
rect 2758 368 2766 371
rect 2770 368 2798 371
rect 2834 368 2918 371
rect 2978 368 3150 371
rect 3350 368 3486 371
rect 3642 368 3646 371
rect 310 362 313 368
rect 42 358 86 361
rect 1198 361 1201 368
rect 2030 362 2033 368
rect 898 358 1462 361
rect 1474 358 1518 361
rect 1546 358 1686 361
rect 1694 358 1830 361
rect 1842 358 1982 361
rect 2010 358 2014 361
rect 2234 358 2246 361
rect 2314 358 2318 361
rect 2378 358 2398 361
rect 2418 358 2462 361
rect 2502 361 2505 368
rect 3214 362 3217 368
rect 3350 362 3353 368
rect 2502 358 2702 361
rect 2738 358 2750 361
rect 2754 358 2766 361
rect 2826 358 2862 361
rect 2938 358 3014 361
rect 3098 358 3150 361
rect 3162 358 3166 361
rect 3218 358 3326 361
rect 3458 358 3462 361
rect 3466 358 3518 361
rect 3522 358 3614 361
rect 3634 358 3638 361
rect 3666 358 3670 361
rect 590 352 593 358
rect 666 348 822 351
rect 830 348 854 351
rect 906 348 974 351
rect 1002 348 1046 351
rect 1050 348 1110 351
rect 1130 348 1142 351
rect 1154 348 1246 351
rect 1398 348 1510 351
rect 1530 348 1550 351
rect 1554 348 1574 351
rect 1694 351 1697 358
rect 2494 352 2497 358
rect 1658 348 1697 351
rect 1802 348 1862 351
rect 1954 348 2030 351
rect 2090 348 2126 351
rect 2330 348 2342 351
rect 2346 348 2350 351
rect 2370 348 2438 351
rect 2474 348 2494 351
rect 2506 348 2566 351
rect 2674 348 2694 351
rect 2722 348 2726 351
rect 2738 348 2750 351
rect 2778 348 2790 351
rect 2850 348 2854 351
rect 2874 348 2878 351
rect 2922 348 2926 351
rect 3018 348 3278 351
rect 3282 348 3358 351
rect 3362 348 3438 351
rect 3482 348 3502 351
rect 3654 351 3657 358
rect 3562 348 3657 351
rect 534 342 537 348
rect 358 338 494 341
rect 554 338 606 341
rect 830 341 833 348
rect 1398 342 1401 348
rect 750 338 833 341
rect 850 338 870 341
rect 906 338 926 341
rect 946 338 1006 341
rect 1018 338 1022 341
rect 1050 338 1105 341
rect 1130 338 1390 341
rect 1426 338 1542 341
rect 1654 338 1662 341
rect 1726 341 1729 348
rect 1666 338 1729 341
rect 1834 338 1838 341
rect 1842 338 1974 341
rect 2034 338 2046 341
rect 2066 338 2073 341
rect 2082 338 2086 341
rect 2238 341 2241 348
rect 2114 338 2241 341
rect 2270 342 2273 348
rect 2286 342 2289 348
rect 2702 342 2705 348
rect 3662 342 3665 348
rect 3758 342 3761 348
rect 2306 338 2334 341
rect 2338 338 2342 341
rect 2418 338 2422 341
rect 2426 338 2462 341
rect 2514 338 2598 341
rect 2714 338 2750 341
rect 2762 338 2790 341
rect 2858 338 2889 341
rect 3066 338 3078 341
rect 3082 338 3137 341
rect 3162 338 3198 341
rect 3226 338 3230 341
rect 3338 338 3382 341
rect 3434 338 3470 341
rect 3578 338 3622 341
rect 3706 338 3710 341
rect 142 332 145 338
rect 358 332 361 338
rect 734 332 737 338
rect 750 332 753 338
rect 1102 332 1105 338
rect 378 328 553 331
rect 550 322 553 328
rect 842 328 934 331
rect 938 328 982 331
rect 1042 328 1094 331
rect 1114 328 1134 331
rect 1234 328 1278 331
rect 1322 328 1382 331
rect 1422 331 1425 338
rect 1742 332 1745 338
rect 1386 328 1425 331
rect 1586 328 1694 331
rect 1866 328 1910 331
rect 1922 328 1958 331
rect 1962 328 1990 331
rect 2026 328 2030 331
rect 2042 328 2054 331
rect 2070 331 2073 338
rect 2070 328 2102 331
rect 2138 328 2230 331
rect 2238 331 2241 338
rect 2886 332 2889 338
rect 3134 332 3137 338
rect 2238 328 2342 331
rect 2386 328 2406 331
rect 2426 328 2534 331
rect 2658 328 2822 331
rect 2826 328 2830 331
rect 2898 328 2958 331
rect 3186 328 3278 331
rect 3302 331 3305 338
rect 3282 328 3297 331
rect 3302 328 3350 331
rect 3378 328 3414 331
rect 3642 328 3822 331
rect 630 321 633 328
rect 630 318 1046 321
rect 1302 321 1305 328
rect 3174 322 3177 328
rect 3294 322 3297 328
rect 3518 322 3521 328
rect 3598 322 3601 328
rect 3622 322 3625 328
rect 1186 318 1305 321
rect 1330 318 1446 321
rect 1482 318 1990 321
rect 1994 318 2214 321
rect 2218 318 2262 321
rect 2266 318 2710 321
rect 2842 318 2854 321
rect 2858 318 2878 321
rect 2894 318 3110 321
rect 3274 318 3278 321
rect 3650 318 3758 321
rect 506 308 518 311
rect 550 311 553 318
rect 710 312 713 318
rect 550 308 582 311
rect 986 308 1070 311
rect 1194 308 1238 311
rect 1242 308 1294 311
rect 1306 308 1334 311
rect 1362 308 1542 311
rect 1554 308 1766 311
rect 1834 308 1870 311
rect 1962 308 2046 311
rect 2050 308 2286 311
rect 2290 308 2542 311
rect 2562 308 2574 311
rect 2894 311 2897 318
rect 2586 308 2897 311
rect 2954 308 3030 311
rect 3114 308 3254 311
rect 3258 308 3286 311
rect 3314 308 3462 311
rect 848 303 850 307
rect 854 303 857 307
rect 862 303 864 307
rect 1880 303 1882 307
rect 1886 303 1889 307
rect 1894 303 1896 307
rect 2904 303 2906 307
rect 2910 303 2913 307
rect 2918 303 2920 307
rect 74 298 86 301
rect 970 298 998 301
rect 1026 298 1214 301
rect 1274 298 1870 301
rect 1926 298 2390 301
rect 2394 298 2470 301
rect 2482 298 2550 301
rect 2570 298 2590 301
rect 2626 298 2678 301
rect 2690 298 2702 301
rect 2810 298 2870 301
rect 2874 298 2894 301
rect 2986 298 2990 301
rect 3154 298 3270 301
rect 3282 298 3406 301
rect 3474 298 3646 301
rect 178 288 286 291
rect 466 288 494 291
rect 922 288 1054 291
rect 1098 288 1254 291
rect 1530 288 1566 291
rect 1578 288 1622 291
rect 1870 291 1873 298
rect 1926 292 1929 298
rect 1634 288 1809 291
rect 1870 288 1926 291
rect 1938 288 1998 291
rect 2046 288 2062 291
rect 2074 288 2118 291
rect 2154 288 2158 291
rect 2226 288 2302 291
rect 2442 288 2446 291
rect 2470 291 2473 298
rect 2470 288 3038 291
rect 3042 288 3318 291
rect 3594 288 3694 291
rect 578 278 598 281
rect 830 281 833 288
rect 818 278 833 281
rect 850 278 950 281
rect 986 278 1014 281
rect 1026 278 1078 281
rect 1098 278 1118 281
rect 1318 281 1321 288
rect 1298 278 1321 281
rect 1502 282 1505 288
rect 1514 278 1518 281
rect 1582 278 1654 281
rect 1658 278 1726 281
rect 1730 278 1798 281
rect 1806 281 1809 288
rect 2030 282 2033 288
rect 2046 282 2049 288
rect 2206 282 2209 288
rect 2214 282 2217 288
rect 1806 278 1974 281
rect 2058 278 2062 281
rect 2066 278 2102 281
rect 2114 278 2118 281
rect 2138 278 2198 281
rect 2234 278 2238 281
rect 2250 278 2310 281
rect 2362 278 2590 281
rect 2874 278 2934 281
rect 2982 278 3014 281
rect 3018 278 3126 281
rect 3274 278 3326 281
rect 3446 281 3449 288
rect 3346 278 3449 281
rect 3506 278 3710 281
rect 70 272 73 278
rect 286 272 289 278
rect 478 272 481 278
rect 550 272 553 278
rect 1534 272 1537 278
rect 1582 272 1585 278
rect 2862 272 2865 278
rect 2982 272 2985 278
rect 3190 272 3193 278
rect 554 268 670 271
rect 762 268 974 271
rect 1042 268 1102 271
rect 1114 268 1174 271
rect 1386 268 1510 271
rect 1514 268 1518 271
rect 1578 268 1582 271
rect 1594 268 1598 271
rect 1618 268 1622 271
rect 1690 268 1750 271
rect 1754 268 1758 271
rect 1762 268 1814 271
rect 1818 268 2014 271
rect 2018 268 2574 271
rect 2594 268 2598 271
rect 2610 268 2846 271
rect 2990 268 3022 271
rect 3206 271 3209 278
rect 3206 268 3246 271
rect 3338 268 3350 271
rect 3506 268 3574 271
rect 186 258 342 261
rect 346 258 422 261
rect 562 258 566 261
rect 570 258 598 261
rect 954 258 966 261
rect 970 258 1014 261
rect 1026 258 1046 261
rect 1090 258 1142 261
rect 1170 258 1182 261
rect 1218 258 1878 261
rect 1882 258 1958 261
rect 1978 258 2614 261
rect 2618 258 2790 261
rect 2842 258 2870 261
rect 2990 261 2993 268
rect 3150 262 3153 268
rect 3614 262 3617 268
rect 2938 258 2993 261
rect 3010 258 3014 261
rect 3154 258 3190 261
rect 3282 258 3286 261
rect 3290 258 3318 261
rect 662 252 665 258
rect 338 248 374 251
rect 986 248 1094 251
rect 1106 248 1182 251
rect 1402 248 1462 251
rect 1466 248 1526 251
rect 1546 248 1614 251
rect 1626 248 1630 251
rect 1642 248 1670 251
rect 1706 248 1710 251
rect 1722 248 1742 251
rect 1762 248 1766 251
rect 1778 248 1782 251
rect 1794 248 1814 251
rect 1930 248 1934 251
rect 1978 248 2094 251
rect 2098 248 2150 251
rect 2154 248 2158 251
rect 2162 248 2166 251
rect 2202 248 2206 251
rect 2242 248 2478 251
rect 2506 248 2510 251
rect 2522 248 2590 251
rect 2846 248 2902 251
rect 3018 248 3022 251
rect 3106 248 3142 251
rect 3302 248 3326 251
rect 3498 248 3710 251
rect 994 238 1030 241
rect 1074 238 1142 241
rect 1178 238 1182 241
rect 1202 238 1438 241
rect 1534 241 1537 248
rect 2846 242 2849 248
rect 1498 238 1537 241
rect 1562 238 1566 241
rect 1618 238 1833 241
rect 1850 238 1878 241
rect 1954 238 1982 241
rect 2002 238 2182 241
rect 2186 238 2190 241
rect 2226 238 2270 241
rect 2274 238 2630 241
rect 2634 238 2662 241
rect 2666 238 2838 241
rect 2942 241 2945 248
rect 2890 238 2945 241
rect 3302 242 3305 248
rect 634 228 750 231
rect 978 228 1806 231
rect 1830 231 1833 238
rect 1830 228 2038 231
rect 2042 228 2078 231
rect 2210 228 2534 231
rect 2650 228 2974 231
rect 2986 228 3126 231
rect 3130 228 3302 231
rect 3306 228 3766 231
rect 226 218 374 221
rect 962 218 998 221
rect 1006 218 1086 221
rect 1218 218 1438 221
rect 1586 218 1638 221
rect 1650 218 1782 221
rect 1986 218 2310 221
rect 2314 218 2470 221
rect 2482 218 2774 221
rect 2778 218 2830 221
rect 2842 218 2878 221
rect 2898 218 3278 221
rect 3282 218 3289 221
rect 3298 218 3534 221
rect 3722 218 3734 221
rect 90 208 110 211
rect 114 208 270 211
rect 1006 211 1009 218
rect 498 208 1009 211
rect 1066 208 1342 211
rect 1438 211 1441 218
rect 1438 208 2006 211
rect 2170 208 2190 211
rect 2234 208 2350 211
rect 2562 208 2870 211
rect 2874 208 3054 211
rect 3058 208 3086 211
rect 3450 208 3454 211
rect 3538 208 3758 211
rect 344 203 346 207
rect 350 203 353 207
rect 358 203 360 207
rect 1360 203 1362 207
rect 1366 203 1369 207
rect 1374 203 1376 207
rect 2014 202 2017 208
rect 2384 203 2386 207
rect 2390 203 2393 207
rect 2398 203 2400 207
rect 3408 203 3410 207
rect 3414 203 3417 207
rect 3422 203 3424 207
rect 594 198 662 201
rect 666 198 1134 201
rect 1138 198 1350 201
rect 1626 198 1734 201
rect 2022 198 2214 201
rect 2274 198 2286 201
rect 2578 198 2910 201
rect 2966 198 3030 201
rect 3066 198 3102 201
rect 3106 198 3310 201
rect 3570 198 3742 201
rect 122 188 158 191
rect 522 188 550 191
rect 754 188 1158 191
rect 1162 188 1454 191
rect 1458 188 1662 191
rect 2022 191 2025 198
rect 1906 188 2025 191
rect 2050 188 2182 191
rect 2186 188 2422 191
rect 2426 188 2430 191
rect 2474 188 2478 191
rect 2634 188 2654 191
rect 2742 188 2814 191
rect 2966 191 2969 198
rect 2818 188 2969 191
rect 2978 188 3006 191
rect 3074 188 3078 191
rect 3410 188 3590 191
rect 2742 182 2745 188
rect 330 178 670 181
rect 986 178 1022 181
rect 1034 178 1070 181
rect 1074 178 1273 181
rect 1282 178 1478 181
rect 1618 178 1654 181
rect 1666 178 1702 181
rect 1922 178 1990 181
rect 1994 178 2718 181
rect 2930 178 2974 181
rect 2978 178 3238 181
rect 3546 178 3582 181
rect 1270 172 1273 178
rect 722 168 806 171
rect 1002 168 1030 171
rect 1050 168 1102 171
rect 1106 168 1118 171
rect 1134 168 1262 171
rect 1290 168 1846 171
rect 1962 168 2118 171
rect 2122 168 2174 171
rect 2282 168 2430 171
rect 2714 168 2958 171
rect 2962 168 3158 171
rect 3554 168 3558 171
rect 3714 168 3718 171
rect 614 161 617 168
rect 354 158 617 161
rect 642 158 766 161
rect 982 161 985 168
rect 1134 162 1137 168
rect 906 158 985 161
rect 1034 158 1054 161
rect 1058 158 1065 161
rect 1194 158 1198 161
rect 1306 158 1566 161
rect 2090 158 2102 161
rect 2106 158 2166 161
rect 2234 158 2238 161
rect 2258 158 2358 161
rect 2402 158 2486 161
rect 2490 158 2518 161
rect 2690 158 2710 161
rect 2714 158 2942 161
rect 2946 158 2998 161
rect 3002 158 3006 161
rect 3042 158 3078 161
rect 3566 161 3569 168
rect 3566 158 3574 161
rect 1214 152 1217 158
rect -26 151 -22 152
rect -26 148 6 151
rect 90 148 166 151
rect 170 148 198 151
rect 602 148 638 151
rect 642 148 694 151
rect 698 148 718 151
rect 994 148 1006 151
rect 1010 148 1054 151
rect 1114 148 1182 151
rect 1234 148 1238 151
rect 1426 148 1518 151
rect 1702 151 1705 158
rect 1690 148 1705 151
rect 1818 148 1926 151
rect 2138 148 2142 151
rect 2162 148 2190 151
rect 2210 148 2278 151
rect 2722 148 2726 151
rect 2834 148 2886 151
rect 2890 148 2894 151
rect 2970 148 2990 151
rect 3010 148 3049 151
rect 3162 148 3166 151
rect 3554 148 3558 151
rect 3598 151 3601 158
rect 3598 148 3606 151
rect 3610 148 3622 151
rect 3662 151 3665 158
rect 3718 152 3721 158
rect 3626 148 3665 151
rect 3682 148 3686 151
rect 38 142 41 148
rect 42 138 262 141
rect 514 138 598 141
rect 610 138 630 141
rect 634 138 686 141
rect 690 138 718 141
rect 970 138 1142 141
rect 1178 138 1206 141
rect 1210 138 1214 141
rect 1218 138 1238 141
rect 1366 141 1369 148
rect 1266 138 1369 141
rect 1982 141 1985 148
rect 2150 142 2153 148
rect 1982 138 2126 141
rect 2186 138 2222 141
rect 2234 138 2238 141
rect 2342 141 2345 148
rect 3046 142 3049 148
rect 3422 142 3425 148
rect 2250 138 2345 141
rect 2690 138 2694 141
rect 2738 138 2846 141
rect 2930 138 2998 141
rect 3002 138 3014 141
rect 3026 138 3030 141
rect 3146 138 3222 141
rect 3290 138 3294 141
rect 3306 138 3366 141
rect 3674 138 3678 141
rect 510 131 513 138
rect 258 128 513 131
rect 818 128 1014 131
rect 1018 128 1070 131
rect 1082 128 1214 131
rect 1382 128 1462 131
rect 1742 131 1745 138
rect 2558 132 2561 138
rect 1466 128 1745 131
rect 1898 128 1918 131
rect 2802 128 2822 131
rect 2826 128 3006 131
rect 3142 131 3145 138
rect 3010 128 3145 131
rect 3406 131 3409 138
rect 3234 128 3409 131
rect 3498 128 3662 131
rect 3706 128 3710 131
rect 1382 122 1385 128
rect 282 118 774 121
rect 782 118 1278 121
rect 2126 121 2129 128
rect 1762 118 2129 121
rect 2678 121 2681 128
rect 2282 118 2681 121
rect 2850 118 3022 121
rect 3098 118 3310 121
rect 3322 118 3574 121
rect 782 111 785 118
rect 138 108 785 111
rect 1258 108 1318 111
rect 2010 108 2206 111
rect 2234 108 2294 111
rect 2374 108 2486 111
rect 2490 108 2646 111
rect 3130 108 3238 111
rect 3362 108 3606 111
rect 3698 108 3742 111
rect 848 103 850 107
rect 854 103 857 107
rect 862 103 864 107
rect 1880 103 1882 107
rect 1886 103 1889 107
rect 1894 103 1896 107
rect 2374 102 2377 108
rect 2904 103 2906 107
rect 2910 103 2913 107
rect 2918 103 2920 107
rect 602 98 710 101
rect 730 98 734 101
rect 890 98 918 101
rect 922 98 1518 101
rect 1522 98 1566 101
rect 1570 98 1790 101
rect 1794 98 1814 101
rect 1818 98 1830 101
rect 2002 98 2294 101
rect 2306 98 2374 101
rect 2610 98 2854 101
rect 3114 98 3134 101
rect 3402 98 3718 101
rect 3142 92 3145 98
rect 490 88 622 91
rect 626 88 734 91
rect 770 88 1118 91
rect 1122 88 1310 91
rect 1314 88 1318 91
rect 1618 88 1646 91
rect 2106 88 2214 91
rect 2506 88 2582 91
rect 2858 88 3094 91
rect 3450 88 3598 91
rect 3634 88 3638 91
rect 3690 88 3734 91
rect 118 81 121 88
rect 118 78 254 81
rect 486 81 489 88
rect 418 78 489 81
rect 906 78 910 81
rect 1530 78 1566 81
rect 1630 78 1750 81
rect 1754 78 1806 81
rect 2094 81 2097 88
rect 3430 82 3433 88
rect 2094 78 2254 81
rect 2294 78 2758 81
rect 3138 78 3142 81
rect 3490 78 3681 81
rect 3714 78 3718 81
rect 502 72 505 78
rect 750 72 753 78
rect 1102 71 1105 78
rect 1630 72 1633 78
rect 1102 68 1118 71
rect 1490 68 1526 71
rect 2078 71 2081 78
rect 2294 72 2297 78
rect 2494 72 2497 78
rect 2670 72 2673 78
rect 2078 68 2102 71
rect 2186 68 2206 71
rect 2210 68 2214 71
rect 2510 68 2606 71
rect 2686 68 2742 71
rect 2886 71 2889 78
rect 2990 71 2993 78
rect 2886 68 2993 71
rect 3050 68 3190 71
rect 3246 71 3249 78
rect 3234 68 3249 71
rect 3334 72 3337 78
rect 3678 72 3681 78
rect 3758 72 3761 78
rect 3354 68 3358 71
rect 3474 68 3550 71
rect 3586 68 3590 71
rect 3682 68 3694 71
rect 2038 62 2041 68
rect 2510 62 2513 68
rect 2686 62 2689 68
rect 3390 62 3393 68
rect 314 58 558 61
rect 578 58 582 61
rect 622 58 630 61
rect 634 58 646 61
rect 962 58 1046 61
rect 1162 58 1246 61
rect 1970 58 2038 61
rect 2138 58 2222 61
rect 2570 58 2630 61
rect 2746 58 2782 61
rect 2834 58 2846 61
rect 2914 58 2950 61
rect 3130 58 3318 61
rect 3370 58 3374 61
rect 3482 58 3486 61
rect 3530 58 3614 61
rect 3658 58 3686 61
rect 3714 58 3766 61
rect -26 51 -22 52
rect -26 48 6 51
rect 242 48 262 51
rect 1698 48 2406 51
rect 2410 48 2854 51
rect 3362 48 3641 51
rect 3650 48 3726 51
rect 3330 38 3334 41
rect 3378 38 3382 41
rect 3394 38 3454 41
rect 3638 41 3641 48
rect 3638 38 3750 41
rect 1346 28 1998 31
rect 2002 28 2014 31
rect 3590 31 3593 38
rect 3346 28 3646 31
rect 1214 12 1217 18
rect 1278 12 1281 18
rect 1926 12 1929 18
rect 2094 12 2097 18
rect 730 8 734 11
rect 770 8 782 11
rect 1090 8 1102 11
rect 1234 8 1254 11
rect 2498 8 2510 11
rect 344 3 346 7
rect 350 3 353 7
rect 358 3 360 7
rect 1360 3 1362 7
rect 1366 3 1369 7
rect 1374 3 1376 7
rect 2384 3 2386 7
rect 2390 3 2393 7
rect 2398 3 2400 7
rect 3408 3 3410 7
rect 3414 3 3417 7
rect 3422 3 3424 7
<< m4contact >>
rect 346 3603 350 3607
rect 354 3603 357 3607
rect 357 3603 358 3607
rect 1362 3603 1366 3607
rect 1370 3603 1373 3607
rect 1373 3603 1374 3607
rect 2386 3603 2390 3607
rect 2394 3603 2397 3607
rect 2397 3603 2398 3607
rect 3410 3603 3414 3607
rect 3418 3603 3421 3607
rect 3421 3603 3422 3607
rect 422 3598 426 3602
rect 894 3598 898 3602
rect 1478 3598 1482 3602
rect 1502 3598 1506 3602
rect 1958 3598 1962 3602
rect 1070 3588 1074 3592
rect 1270 3588 1274 3592
rect 1334 3588 1338 3592
rect 1574 3588 1578 3592
rect 1606 3588 1610 3592
rect 1758 3588 1762 3592
rect 1798 3588 1802 3592
rect 1902 3588 1906 3592
rect 2070 3588 2074 3592
rect 2230 3588 2234 3592
rect 2406 3588 2410 3592
rect 2974 3588 2978 3592
rect 3334 3588 3338 3592
rect 1398 3578 1402 3582
rect 2070 3568 2074 3572
rect 3534 3568 3538 3572
rect 1862 3558 1866 3562
rect 2126 3558 2130 3562
rect 734 3548 738 3552
rect 3150 3548 3154 3552
rect 3334 3548 3338 3552
rect 3614 3548 3618 3552
rect 3662 3548 3666 3552
rect 670 3538 674 3542
rect 902 3538 906 3542
rect 1062 3538 1066 3542
rect 1582 3538 1586 3542
rect 1662 3538 1666 3542
rect 1798 3538 1802 3542
rect 2006 3538 2010 3542
rect 2166 3538 2170 3542
rect 2398 3538 2402 3542
rect 2574 3538 2578 3542
rect 3206 3538 3210 3542
rect 3326 3538 3330 3542
rect 3654 3538 3658 3542
rect 3734 3538 3738 3542
rect 966 3528 970 3532
rect 1302 3528 1306 3532
rect 1974 3528 1978 3532
rect 1982 3528 1986 3532
rect 2278 3528 2282 3532
rect 2486 3528 2490 3532
rect 3150 3528 3154 3532
rect 3262 3528 3266 3532
rect 3598 3528 3602 3532
rect 3710 3528 3714 3532
rect 3726 3528 3730 3532
rect 294 3518 298 3522
rect 1286 3518 1290 3522
rect 2926 3518 2930 3522
rect 2942 3518 2946 3522
rect 3558 3518 3562 3522
rect 430 3508 434 3512
rect 870 3508 874 3512
rect 1142 3508 1146 3512
rect 2238 3508 2242 3512
rect 2270 3508 2274 3512
rect 2870 3508 2874 3512
rect 3254 3508 3258 3512
rect 850 3503 854 3507
rect 858 3503 861 3507
rect 861 3503 862 3507
rect 1882 3503 1886 3507
rect 1890 3503 1893 3507
rect 1893 3503 1894 3507
rect 2906 3503 2910 3507
rect 2914 3503 2917 3507
rect 2917 3503 2918 3507
rect 1286 3498 1290 3502
rect 2926 3498 2930 3502
rect 3598 3488 3602 3492
rect 3606 3488 3610 3492
rect 678 3478 682 3482
rect 1878 3478 1882 3482
rect 2894 3478 2898 3482
rect 3566 3478 3570 3482
rect 3582 3478 3586 3482
rect 3718 3478 3722 3482
rect 702 3468 706 3472
rect 894 3468 898 3472
rect 1422 3468 1426 3472
rect 2022 3468 2026 3472
rect 2574 3468 2578 3472
rect 3510 3468 3514 3472
rect 3630 3468 3634 3472
rect 3742 3468 3746 3472
rect 6 3458 10 3462
rect 198 3458 202 3462
rect 2126 3458 2130 3462
rect 2262 3458 2266 3462
rect 2550 3458 2554 3462
rect 3686 3458 3690 3462
rect 3702 3458 3706 3462
rect 1750 3448 1754 3452
rect 2558 3448 2562 3452
rect 2958 3448 2962 3452
rect 3014 3448 3018 3452
rect 3190 3448 3194 3452
rect 3206 3448 3210 3452
rect 3638 3448 3642 3452
rect 3774 3448 3778 3452
rect 558 3438 562 3442
rect 2334 3438 2338 3442
rect 3262 3438 3266 3442
rect 3534 3438 3538 3442
rect 3590 3438 3594 3442
rect 3614 3438 3618 3442
rect 3654 3438 3658 3442
rect 582 3428 586 3432
rect 870 3428 874 3432
rect 2558 3428 2562 3432
rect 3670 3428 3674 3432
rect 942 3418 946 3422
rect 1070 3418 1074 3422
rect 1606 3418 1610 3422
rect 1870 3418 1874 3422
rect 2222 3418 2226 3422
rect 2414 3418 2418 3422
rect 3262 3418 3266 3422
rect 3278 3418 3282 3422
rect 3670 3418 3674 3422
rect 734 3408 738 3412
rect 1318 3408 1322 3412
rect 1382 3408 1386 3412
rect 2374 3408 2378 3412
rect 3286 3408 3290 3412
rect 3294 3408 3298 3412
rect 3542 3408 3546 3412
rect 346 3403 350 3407
rect 354 3403 357 3407
rect 357 3403 358 3407
rect 1362 3403 1366 3407
rect 1370 3403 1373 3407
rect 1373 3403 1374 3407
rect 2386 3403 2390 3407
rect 2394 3403 2397 3407
rect 2397 3403 2398 3407
rect 3410 3403 3414 3407
rect 3418 3403 3421 3407
rect 3421 3403 3422 3407
rect 558 3398 562 3402
rect 1574 3398 1578 3402
rect 1750 3398 1754 3402
rect 1798 3398 1802 3402
rect 3374 3398 3378 3402
rect 238 3388 242 3392
rect 2278 3388 2282 3392
rect 3198 3388 3202 3392
rect 3342 3388 3346 3392
rect 3678 3388 3682 3392
rect 1302 3378 1306 3382
rect 3014 3378 3018 3382
rect 3182 3378 3186 3382
rect 3270 3378 3274 3382
rect 3374 3378 3378 3382
rect 3726 3378 3730 3382
rect 1310 3368 1314 3372
rect 1318 3368 1322 3372
rect 1654 3368 1658 3372
rect 2550 3368 2554 3372
rect 3342 3368 3346 3372
rect 1262 3358 1266 3362
rect 2406 3358 2410 3362
rect 2894 3358 2898 3362
rect 3022 3358 3026 3362
rect 3414 3358 3418 3362
rect 3518 3358 3522 3362
rect 3694 3358 3698 3362
rect 1926 3348 1930 3352
rect 2318 3348 2322 3352
rect 3286 3348 3290 3352
rect 3646 3348 3650 3352
rect 774 3338 778 3342
rect 982 3338 986 3342
rect 1110 3338 1114 3342
rect 1358 3338 1362 3342
rect 1846 3338 1850 3342
rect 2110 3338 2114 3342
rect 2166 3338 2170 3342
rect 3678 3338 3682 3342
rect 3718 3338 3722 3342
rect 678 3328 682 3332
rect 950 3328 954 3332
rect 1318 3328 1322 3332
rect 2198 3328 2202 3332
rect 2302 3328 2306 3332
rect 2926 3328 2930 3332
rect 3174 3328 3178 3332
rect 502 3318 506 3322
rect 1182 3318 1186 3322
rect 1382 3318 1386 3322
rect 1398 3318 1402 3322
rect 2126 3318 2130 3322
rect 2246 3318 2250 3322
rect 2302 3318 2306 3322
rect 2358 3318 2362 3322
rect 3006 3318 3010 3322
rect 3270 3318 3274 3322
rect 3278 3318 3282 3322
rect 3622 3318 3626 3322
rect 3758 3318 3762 3322
rect 1862 3308 1866 3312
rect 2022 3308 2026 3312
rect 2670 3308 2674 3312
rect 850 3303 854 3307
rect 858 3303 861 3307
rect 861 3303 862 3307
rect 1882 3303 1886 3307
rect 1890 3303 1893 3307
rect 1893 3303 1894 3307
rect 2906 3303 2910 3307
rect 2914 3303 2917 3307
rect 2917 3303 2918 3307
rect 230 3298 234 3302
rect 1022 3298 1026 3302
rect 1134 3298 1138 3302
rect 2014 3298 2018 3302
rect 2926 3298 2930 3302
rect 1326 3288 1330 3292
rect 1414 3288 1418 3292
rect 1510 3288 1514 3292
rect 3038 3288 3042 3292
rect 942 3278 946 3282
rect 950 3278 954 3282
rect 1782 3278 1786 3282
rect 2870 3278 2874 3282
rect 3006 3278 3010 3282
rect 3174 3278 3178 3282
rect 3550 3278 3554 3282
rect 134 3268 138 3272
rect 286 3268 290 3272
rect 782 3268 786 3272
rect 1158 3268 1162 3272
rect 1654 3268 1658 3272
rect 1806 3268 1810 3272
rect 2902 3268 2906 3272
rect 2966 3268 2970 3272
rect 3006 3268 3010 3272
rect 3062 3268 3066 3272
rect 3174 3268 3178 3272
rect 3766 3268 3770 3272
rect 454 3258 458 3262
rect 606 3258 610 3262
rect 1294 3258 1298 3262
rect 1398 3258 1402 3262
rect 2550 3258 2554 3262
rect 3014 3258 3018 3262
rect 3318 3258 3322 3262
rect 3374 3258 3378 3262
rect 3542 3258 3546 3262
rect 3694 3258 3698 3262
rect 318 3248 322 3252
rect 510 3248 514 3252
rect 558 3248 562 3252
rect 590 3248 594 3252
rect 766 3248 770 3252
rect 1094 3248 1098 3252
rect 1302 3248 1306 3252
rect 1894 3248 1898 3252
rect 2886 3248 2890 3252
rect 3150 3248 3154 3252
rect 3550 3248 3554 3252
rect 110 3238 114 3242
rect 742 3238 746 3242
rect 1262 3238 1266 3242
rect 1270 3238 1274 3242
rect 1310 3238 1314 3242
rect 1406 3238 1410 3242
rect 2166 3238 2170 3242
rect 3534 3238 3538 3242
rect 1286 3228 1290 3232
rect 1750 3228 1754 3232
rect 2190 3228 2194 3232
rect 3718 3228 3722 3232
rect 966 3218 970 3222
rect 1798 3208 1802 3212
rect 346 3203 350 3207
rect 354 3203 357 3207
rect 357 3203 358 3207
rect 1362 3203 1366 3207
rect 1370 3203 1373 3207
rect 1373 3203 1374 3207
rect 2386 3203 2390 3207
rect 2394 3203 2397 3207
rect 2397 3203 2398 3207
rect 3410 3203 3414 3207
rect 3418 3203 3421 3207
rect 3421 3203 3422 3207
rect 1710 3198 1714 3202
rect 1934 3198 1938 3202
rect 2062 3198 2066 3202
rect 2310 3198 2314 3202
rect 318 3188 322 3192
rect 1318 3188 1322 3192
rect 3286 3188 3290 3192
rect 3590 3188 3594 3192
rect 574 3178 578 3182
rect 886 3178 890 3182
rect 1350 3178 1354 3182
rect 2670 3178 2674 3182
rect 974 3168 978 3172
rect 1790 3168 1794 3172
rect 2630 3168 2634 3172
rect 3158 3168 3162 3172
rect 726 3158 730 3162
rect 998 3158 1002 3162
rect 1262 3158 1266 3162
rect 1526 3158 1530 3162
rect 1798 3158 1802 3162
rect 1910 3158 1914 3162
rect 2078 3158 2082 3162
rect 2150 3158 2154 3162
rect 2230 3158 2234 3162
rect 2590 3158 2594 3162
rect 3134 3158 3138 3162
rect 3350 3158 3354 3162
rect 3526 3158 3530 3162
rect 3622 3158 3626 3162
rect 814 3148 818 3152
rect 1854 3148 1858 3152
rect 2022 3148 2026 3152
rect 2254 3148 2258 3152
rect 2294 3148 2298 3152
rect 6 3138 10 3142
rect 726 3138 730 3142
rect 942 3138 946 3142
rect 974 3138 978 3142
rect 1934 3138 1938 3142
rect 2302 3138 2306 3142
rect 2518 3138 2522 3142
rect 2598 3138 2602 3142
rect 502 3128 506 3132
rect 598 3128 602 3132
rect 758 3128 762 3132
rect 1966 3128 1970 3132
rect 2038 3128 2042 3132
rect 2238 3128 2242 3132
rect 2326 3128 2330 3132
rect 2470 3128 2474 3132
rect 2774 3128 2778 3132
rect 3030 3128 3034 3132
rect 758 3118 762 3122
rect 950 3118 954 3122
rect 1542 3118 1546 3122
rect 1742 3118 1746 3122
rect 1758 3118 1762 3122
rect 2118 3118 2122 3122
rect 2454 3118 2458 3122
rect 2590 3118 2594 3122
rect 2678 3118 2682 3122
rect 574 3108 578 3112
rect 1094 3108 1098 3112
rect 1470 3108 1474 3112
rect 1614 3108 1618 3112
rect 1678 3108 1682 3112
rect 2222 3108 2226 3112
rect 3118 3108 3122 3112
rect 3198 3108 3202 3112
rect 850 3103 854 3107
rect 858 3103 861 3107
rect 861 3103 862 3107
rect 1882 3103 1886 3107
rect 1890 3103 1893 3107
rect 1893 3103 1894 3107
rect 2906 3103 2910 3107
rect 2914 3103 2917 3107
rect 2917 3103 2918 3107
rect 1406 3098 1410 3102
rect 1710 3098 1714 3102
rect 1870 3098 1874 3102
rect 2126 3098 2130 3102
rect 2246 3098 2250 3102
rect 2286 3098 2290 3102
rect 3302 3098 3306 3102
rect 2030 3088 2034 3092
rect 2278 3088 2282 3092
rect 2806 3088 2810 3092
rect 3694 3088 3698 3092
rect 3750 3088 3754 3092
rect 582 3078 586 3082
rect 782 3078 786 3082
rect 966 3078 970 3082
rect 1654 3078 1658 3082
rect 2006 3078 2010 3082
rect 2574 3078 2578 3082
rect 3182 3078 3186 3082
rect 3534 3078 3538 3082
rect 3614 3078 3618 3082
rect 3710 3078 3714 3082
rect 230 3068 234 3072
rect 566 3068 570 3072
rect 646 3068 650 3072
rect 742 3068 746 3072
rect 1094 3068 1098 3072
rect 1398 3068 1402 3072
rect 1406 3068 1410 3072
rect 1486 3068 1490 3072
rect 1678 3068 1682 3072
rect 1686 3068 1690 3072
rect 1926 3068 1930 3072
rect 2022 3068 2026 3072
rect 2254 3068 2258 3072
rect 2582 3068 2586 3072
rect 3014 3068 3018 3072
rect 3310 3068 3314 3072
rect 3510 3068 3514 3072
rect 222 3058 226 3062
rect 238 3058 242 3062
rect 1422 3058 1426 3062
rect 1550 3058 1554 3062
rect 1998 3058 2002 3062
rect 2134 3058 2138 3062
rect 2158 3058 2162 3062
rect 2262 3058 2266 3062
rect 2270 3058 2274 3062
rect 2302 3058 2306 3062
rect 2438 3058 2442 3062
rect 2462 3058 2466 3062
rect 2614 3058 2618 3062
rect 3062 3058 3066 3062
rect 3206 3058 3210 3062
rect 3622 3058 3626 3062
rect 1238 3048 1242 3052
rect 1598 3048 1602 3052
rect 1670 3048 1674 3052
rect 2006 3048 2010 3052
rect 2422 3048 2426 3052
rect 2694 3048 2698 3052
rect 3118 3048 3122 3052
rect 598 3038 602 3042
rect 662 3038 666 3042
rect 926 3038 930 3042
rect 950 3038 954 3042
rect 1174 3038 1178 3042
rect 1622 3038 1626 3042
rect 1678 3038 1682 3042
rect 1790 3038 1794 3042
rect 2102 3038 2106 3042
rect 2118 3038 2122 3042
rect 2254 3038 2258 3042
rect 2598 3038 2602 3042
rect 2654 3038 2658 3042
rect 3534 3048 3538 3052
rect 3590 3048 3594 3052
rect 3598 3048 3602 3052
rect 3750 3048 3754 3052
rect 3406 3038 3410 3042
rect 3534 3038 3538 3042
rect 366 3028 370 3032
rect 1118 3028 1122 3032
rect 1406 3028 1410 3032
rect 1926 3028 1930 3032
rect 2110 3028 2114 3032
rect 2278 3028 2282 3032
rect 3286 3028 3290 3032
rect 1430 3018 1434 3022
rect 1846 3018 1850 3022
rect 1998 3018 2002 3022
rect 2526 3018 2530 3022
rect 3030 3018 3034 3022
rect 582 3008 586 3012
rect 1518 3008 1522 3012
rect 3142 3008 3146 3012
rect 3558 3008 3562 3012
rect 346 3003 350 3007
rect 354 3003 357 3007
rect 357 3003 358 3007
rect 1362 3003 1366 3007
rect 1370 3003 1373 3007
rect 1373 3003 1374 3007
rect 2386 3003 2390 3007
rect 2394 3003 2397 3007
rect 2397 3003 2398 3007
rect 3410 3003 3414 3007
rect 3418 3003 3421 3007
rect 3421 3003 3422 3007
rect 766 2998 770 3002
rect 894 2998 898 3002
rect 950 2998 954 3002
rect 1390 2998 1394 3002
rect 1878 2998 1882 3002
rect 2126 2998 2130 3002
rect 2582 2998 2586 3002
rect 590 2988 594 2992
rect 918 2988 922 2992
rect 1262 2988 1266 2992
rect 1566 2988 1570 2992
rect 2238 2988 2242 2992
rect 2318 2988 2322 2992
rect 3270 2988 3274 2992
rect 1254 2978 1258 2982
rect 1270 2978 1274 2982
rect 1326 2978 1330 2982
rect 1662 2978 1666 2982
rect 1974 2978 1978 2982
rect 2030 2978 2034 2982
rect 2046 2978 2050 2982
rect 2070 2978 2074 2982
rect 2102 2978 2106 2982
rect 2614 2978 2618 2982
rect 3126 2978 3130 2982
rect 3342 2978 3346 2982
rect 710 2968 714 2972
rect 1046 2968 1050 2972
rect 1230 2968 1234 2972
rect 1550 2968 1554 2972
rect 1606 2968 1610 2972
rect 1686 2968 1690 2972
rect 2006 2968 2010 2972
rect 2054 2968 2058 2972
rect 2190 2968 2194 2972
rect 2222 2968 2226 2972
rect 2454 2968 2458 2972
rect 2550 2968 2554 2972
rect 3510 2968 3514 2972
rect 910 2958 914 2962
rect 926 2958 930 2962
rect 1270 2958 1274 2962
rect 1286 2958 1290 2962
rect 1326 2958 1330 2962
rect 1478 2958 1482 2962
rect 1726 2958 1730 2962
rect 2974 2958 2978 2962
rect 3158 2958 3162 2962
rect 3318 2958 3322 2962
rect 3390 2958 3394 2962
rect 3494 2958 3498 2962
rect 3654 2958 3658 2962
rect 614 2948 618 2952
rect 838 2948 842 2952
rect 942 2948 946 2952
rect 1942 2948 1946 2952
rect 2462 2948 2466 2952
rect 3334 2948 3338 2952
rect 3382 2948 3386 2952
rect 3462 2948 3466 2952
rect 3622 2948 3626 2952
rect 3678 2948 3682 2952
rect 318 2938 322 2942
rect 550 2938 554 2942
rect 942 2938 946 2942
rect 1238 2938 1242 2942
rect 1270 2938 1274 2942
rect 1446 2938 1450 2942
rect 1510 2938 1514 2942
rect 1526 2938 1530 2942
rect 1542 2938 1546 2942
rect 1598 2938 1602 2942
rect 1614 2938 1618 2942
rect 2006 2938 2010 2942
rect 2062 2938 2066 2942
rect 2070 2938 2074 2942
rect 2134 2938 2138 2942
rect 2502 2938 2506 2942
rect 2710 2938 2714 2942
rect 3174 2938 3178 2942
rect 3302 2938 3306 2942
rect 3510 2938 3514 2942
rect 3694 2938 3698 2942
rect 574 2928 578 2932
rect 694 2928 698 2932
rect 750 2928 754 2932
rect 758 2928 762 2932
rect 974 2928 978 2932
rect 1302 2928 1306 2932
rect 1406 2928 1410 2932
rect 1622 2928 1626 2932
rect 1830 2928 1834 2932
rect 1846 2928 1850 2932
rect 2014 2928 2018 2932
rect 2142 2928 2146 2932
rect 2206 2928 2210 2932
rect 2342 2928 2346 2932
rect 2374 2928 2378 2932
rect 2470 2928 2474 2932
rect 2606 2928 2610 2932
rect 2662 2928 2666 2932
rect 2774 2928 2778 2932
rect 3550 2928 3554 2932
rect 3758 2928 3762 2932
rect 886 2918 890 2922
rect 1510 2918 1514 2922
rect 1662 2918 1666 2922
rect 1862 2918 1866 2922
rect 1878 2918 1882 2922
rect 2270 2918 2274 2922
rect 2310 2918 2314 2922
rect 2926 2918 2930 2922
rect 3670 2918 3674 2922
rect 1518 2908 1522 2912
rect 1870 2908 1874 2912
rect 1902 2908 1906 2912
rect 2118 2908 2122 2912
rect 2318 2908 2322 2912
rect 2486 2908 2490 2912
rect 2878 2908 2882 2912
rect 850 2903 854 2907
rect 858 2903 861 2907
rect 861 2903 862 2907
rect 1882 2903 1886 2907
rect 1890 2903 1893 2907
rect 1893 2903 1894 2907
rect 2906 2903 2910 2907
rect 2914 2903 2917 2907
rect 2917 2903 2918 2907
rect 334 2898 338 2902
rect 782 2898 786 2902
rect 1678 2898 1682 2902
rect 1694 2898 1698 2902
rect 2046 2898 2050 2902
rect 2726 2898 2730 2902
rect 3278 2898 3282 2902
rect 3294 2898 3298 2902
rect 982 2888 986 2892
rect 1182 2888 1186 2892
rect 2198 2888 2202 2892
rect 2886 2888 2890 2892
rect 3198 2888 3202 2892
rect 3206 2888 3210 2892
rect 3486 2888 3490 2892
rect 3750 2888 3754 2892
rect 230 2878 234 2882
rect 1478 2878 1482 2882
rect 1502 2878 1506 2882
rect 1798 2878 1802 2882
rect 1870 2878 1874 2882
rect 2094 2878 2098 2882
rect 2286 2878 2290 2882
rect 2694 2878 2698 2882
rect 2806 2878 2810 2882
rect 2822 2878 2826 2882
rect 2830 2878 2834 2882
rect 2926 2878 2930 2882
rect 3542 2878 3546 2882
rect 3654 2878 3658 2882
rect 3702 2878 3706 2882
rect 454 2868 458 2872
rect 814 2868 818 2872
rect 862 2868 866 2872
rect 1094 2868 1098 2872
rect 1206 2868 1210 2872
rect 1294 2868 1298 2872
rect 1302 2868 1306 2872
rect 1478 2868 1482 2872
rect 1702 2868 1706 2872
rect 1782 2868 1786 2872
rect 2014 2868 2018 2872
rect 2022 2868 2026 2872
rect 2334 2868 2338 2872
rect 2350 2868 2354 2872
rect 2470 2868 2474 2872
rect 2622 2868 2626 2872
rect 3566 2868 3570 2872
rect 3622 2868 3626 2872
rect 38 2858 42 2862
rect 62 2858 66 2862
rect 758 2858 762 2862
rect 1070 2858 1074 2862
rect 1182 2858 1186 2862
rect 1558 2858 1562 2862
rect 1902 2858 1906 2862
rect 2062 2858 2066 2862
rect 2078 2858 2082 2862
rect 2142 2858 2146 2862
rect 2166 2858 2170 2862
rect 2214 2858 2218 2862
rect 2222 2858 2226 2862
rect 2278 2858 2282 2862
rect 2302 2858 2306 2862
rect 2390 2858 2394 2862
rect 2438 2858 2442 2862
rect 2582 2858 2586 2862
rect 2638 2858 2642 2862
rect 2710 2858 2714 2862
rect 3438 2858 3442 2862
rect 3726 2858 3730 2862
rect 126 2848 130 2852
rect 246 2848 250 2852
rect 1198 2848 1202 2852
rect 1350 2848 1354 2852
rect 1606 2848 1610 2852
rect 1638 2848 1642 2852
rect 2310 2848 2314 2852
rect 2358 2848 2362 2852
rect 2550 2848 2554 2852
rect 2654 2848 2658 2852
rect 2662 2848 2666 2852
rect 2694 2848 2698 2852
rect 2726 2848 2730 2852
rect 3046 2848 3050 2852
rect 3350 2848 3354 2852
rect 3390 2848 3394 2852
rect 110 2838 114 2842
rect 566 2838 570 2842
rect 710 2838 714 2842
rect 870 2838 874 2842
rect 1046 2838 1050 2842
rect 1078 2838 1082 2842
rect 1758 2838 1762 2842
rect 2334 2838 2338 2842
rect 2598 2838 2602 2842
rect 1574 2828 1578 2832
rect 3414 2828 3418 2832
rect 894 2818 898 2822
rect 2150 2818 2154 2822
rect 2222 2818 2226 2822
rect 686 2808 690 2812
rect 1014 2808 1018 2812
rect 1350 2808 1354 2812
rect 1742 2808 1746 2812
rect 1766 2808 1770 2812
rect 2094 2808 2098 2812
rect 2142 2808 2146 2812
rect 2254 2808 2258 2812
rect 2462 2808 2466 2812
rect 2862 2808 2866 2812
rect 3742 2808 3746 2812
rect 346 2803 350 2807
rect 354 2803 357 2807
rect 357 2803 358 2807
rect 1362 2803 1366 2807
rect 1370 2803 1373 2807
rect 1373 2803 1374 2807
rect 2386 2803 2390 2807
rect 2394 2803 2397 2807
rect 2397 2803 2398 2807
rect 3410 2803 3414 2807
rect 3418 2803 3421 2807
rect 3421 2803 3422 2807
rect 214 2798 218 2802
rect 654 2798 658 2802
rect 2374 2798 2378 2802
rect 2686 2798 2690 2802
rect 886 2788 890 2792
rect 1134 2788 1138 2792
rect 1150 2788 1154 2792
rect 1790 2788 1794 2792
rect 2118 2788 2122 2792
rect 2254 2788 2258 2792
rect 2630 2788 2634 2792
rect 2910 2788 2914 2792
rect 3446 2788 3450 2792
rect 710 2778 714 2782
rect 806 2778 810 2782
rect 1526 2778 1530 2782
rect 2166 2778 2170 2782
rect 3238 2778 3242 2782
rect 550 2768 554 2772
rect 766 2768 770 2772
rect 782 2768 786 2772
rect 1334 2768 1338 2772
rect 1422 2768 1426 2772
rect 2350 2768 2354 2772
rect 2558 2768 2562 2772
rect 2718 2768 2722 2772
rect 2798 2768 2802 2772
rect 3086 2768 3090 2772
rect 3198 2768 3202 2772
rect 3518 2768 3522 2772
rect 3558 2768 3562 2772
rect 3742 2768 3746 2772
rect 614 2758 618 2762
rect 1006 2758 1010 2762
rect 1054 2758 1058 2762
rect 1062 2758 1066 2762
rect 1246 2758 1250 2762
rect 1398 2758 1402 2762
rect 1622 2758 1626 2762
rect 1702 2758 1706 2762
rect 1734 2758 1738 2762
rect 1990 2758 1994 2762
rect 2286 2758 2290 2762
rect 2454 2758 2458 2762
rect 2614 2758 2618 2762
rect 3174 2758 3178 2762
rect 334 2748 338 2752
rect 918 2748 922 2752
rect 1438 2748 1442 2752
rect 1742 2748 1746 2752
rect 1814 2748 1818 2752
rect 1870 2748 1874 2752
rect 1990 2748 1994 2752
rect 2014 2748 2018 2752
rect 2358 2748 2362 2752
rect 2374 2748 2378 2752
rect 2670 2748 2674 2752
rect 3270 2748 3274 2752
rect 3654 2748 3658 2752
rect 134 2738 138 2742
rect 566 2738 570 2742
rect 638 2738 642 2742
rect 822 2738 826 2742
rect 846 2738 850 2742
rect 902 2738 906 2742
rect 958 2738 962 2742
rect 1230 2738 1234 2742
rect 1342 2738 1346 2742
rect 1454 2738 1458 2742
rect 1686 2738 1690 2742
rect 1742 2738 1746 2742
rect 2022 2738 2026 2742
rect 2030 2738 2034 2742
rect 2246 2738 2250 2742
rect 2470 2738 2474 2742
rect 2798 2738 2802 2742
rect 3502 2738 3506 2742
rect 3614 2738 3618 2742
rect 670 2728 674 2732
rect 878 2728 882 2732
rect 934 2728 938 2732
rect 1014 2728 1018 2732
rect 1214 2728 1218 2732
rect 1438 2728 1442 2732
rect 1646 2728 1650 2732
rect 1670 2728 1674 2732
rect 1958 2728 1962 2732
rect 2478 2728 2482 2732
rect 2926 2728 2930 2732
rect 3534 2728 3538 2732
rect 3574 2728 3578 2732
rect 1590 2718 1594 2722
rect 1734 2718 1738 2722
rect 1854 2718 1858 2722
rect 1982 2718 1986 2722
rect 2038 2718 2042 2722
rect 2406 2718 2410 2722
rect 2814 2718 2818 2722
rect 3278 2718 3282 2722
rect 3518 2718 3522 2722
rect 3526 2718 3530 2722
rect 3646 2718 3650 2722
rect 3718 2718 3722 2722
rect 3734 2718 3738 2722
rect 518 2708 522 2712
rect 838 2708 842 2712
rect 894 2708 898 2712
rect 1038 2708 1042 2712
rect 1702 2708 1706 2712
rect 1718 2708 1722 2712
rect 2110 2708 2114 2712
rect 2142 2708 2146 2712
rect 2206 2708 2210 2712
rect 2398 2708 2402 2712
rect 2414 2708 2418 2712
rect 2494 2708 2498 2712
rect 2774 2708 2778 2712
rect 3286 2708 3290 2712
rect 3374 2708 3378 2712
rect 3398 2708 3402 2712
rect 850 2703 854 2707
rect 858 2703 861 2707
rect 861 2703 862 2707
rect 1882 2703 1886 2707
rect 1890 2703 1893 2707
rect 1893 2703 1894 2707
rect 2906 2703 2910 2707
rect 2914 2703 2917 2707
rect 2917 2703 2918 2707
rect 894 2698 898 2702
rect 1494 2698 1498 2702
rect 1870 2698 1874 2702
rect 2446 2698 2450 2702
rect 2694 2698 2698 2702
rect 2702 2698 2706 2702
rect 2854 2698 2858 2702
rect 3526 2698 3530 2702
rect 3558 2698 3562 2702
rect 598 2688 602 2692
rect 606 2688 610 2692
rect 870 2688 874 2692
rect 878 2688 882 2692
rect 1126 2688 1130 2692
rect 1142 2688 1146 2692
rect 1478 2688 1482 2692
rect 1662 2688 1666 2692
rect 2078 2688 2082 2692
rect 2246 2688 2250 2692
rect 2422 2688 2426 2692
rect 2934 2688 2938 2692
rect 3542 2688 3546 2692
rect 3622 2688 3626 2692
rect 758 2678 762 2682
rect 806 2678 810 2682
rect 982 2678 986 2682
rect 1086 2678 1090 2682
rect 1990 2678 1994 2682
rect 2270 2678 2274 2682
rect 2366 2678 2370 2682
rect 2646 2678 2650 2682
rect 2718 2678 2722 2682
rect 3046 2678 3050 2682
rect 3118 2678 3122 2682
rect 3190 2678 3194 2682
rect 630 2668 634 2672
rect 646 2668 650 2672
rect 734 2668 738 2672
rect 1014 2668 1018 2672
rect 1078 2668 1082 2672
rect 1590 2668 1594 2672
rect 1838 2668 1842 2672
rect 2118 2668 2122 2672
rect 2158 2668 2162 2672
rect 2254 2668 2258 2672
rect 2686 2668 2690 2672
rect 2694 2668 2698 2672
rect 2734 2668 2738 2672
rect 2838 2668 2842 2672
rect 2846 2668 2850 2672
rect 2862 2668 2866 2672
rect 2894 2668 2898 2672
rect 3510 2668 3514 2672
rect 334 2658 338 2662
rect 462 2658 466 2662
rect 502 2658 506 2662
rect 942 2658 946 2662
rect 974 2658 978 2662
rect 1038 2658 1042 2662
rect 1246 2658 1250 2662
rect 1766 2658 1770 2662
rect 1806 2658 1810 2662
rect 1822 2658 1826 2662
rect 1830 2658 1834 2662
rect 2150 2658 2154 2662
rect 2726 2658 2730 2662
rect 3182 2658 3186 2662
rect 3214 2658 3218 2662
rect 374 2648 378 2652
rect 582 2648 586 2652
rect 878 2648 882 2652
rect 1198 2648 1202 2652
rect 1726 2648 1730 2652
rect 2278 2648 2282 2652
rect 2406 2648 2410 2652
rect 2422 2648 2426 2652
rect 2862 2648 2866 2652
rect 3078 2648 3082 2652
rect 3550 2648 3554 2652
rect 3774 2648 3778 2652
rect 470 2638 474 2642
rect 718 2638 722 2642
rect 734 2638 738 2642
rect 774 2638 778 2642
rect 2214 2638 2218 2642
rect 2294 2638 2298 2642
rect 2654 2638 2658 2642
rect 2750 2638 2754 2642
rect 2830 2638 2834 2642
rect 2838 2638 2842 2642
rect 2902 2638 2906 2642
rect 3062 2638 3066 2642
rect 3246 2638 3250 2642
rect 3654 2638 3658 2642
rect 846 2628 850 2632
rect 918 2628 922 2632
rect 990 2628 994 2632
rect 1254 2628 1258 2632
rect 1750 2628 1754 2632
rect 1934 2628 1938 2632
rect 1958 2628 1962 2632
rect 2742 2628 2746 2632
rect 982 2618 986 2622
rect 1006 2618 1010 2622
rect 1286 2618 1290 2622
rect 1582 2618 1586 2622
rect 1606 2618 1610 2622
rect 2790 2618 2794 2622
rect 3102 2618 3106 2622
rect 3262 2618 3266 2622
rect 1046 2608 1050 2612
rect 1662 2608 1666 2612
rect 1894 2608 1898 2612
rect 2206 2608 2210 2612
rect 2278 2608 2282 2612
rect 2406 2608 2410 2612
rect 3598 2608 3602 2612
rect 346 2603 350 2607
rect 354 2603 357 2607
rect 357 2603 358 2607
rect 1362 2603 1366 2607
rect 1370 2603 1373 2607
rect 1373 2603 1374 2607
rect 2386 2603 2390 2607
rect 2394 2603 2397 2607
rect 2397 2603 2398 2607
rect 598 2598 602 2602
rect 894 2598 898 2602
rect 2158 2598 2162 2602
rect 2550 2598 2554 2602
rect 2670 2598 2674 2602
rect 3410 2603 3414 2607
rect 3418 2603 3421 2607
rect 3421 2603 3422 2607
rect 3398 2598 3402 2602
rect 3494 2598 3498 2602
rect 798 2588 802 2592
rect 926 2588 930 2592
rect 2294 2588 2298 2592
rect 2710 2588 2714 2592
rect 142 2578 146 2582
rect 958 2578 962 2582
rect 1150 2578 1154 2582
rect 1950 2578 1954 2582
rect 2246 2578 2250 2582
rect 2462 2578 2466 2582
rect 2598 2578 2602 2582
rect 2790 2578 2794 2582
rect 2894 2578 2898 2582
rect 3414 2578 3418 2582
rect 3590 2578 3594 2582
rect 766 2568 770 2572
rect 894 2568 898 2572
rect 950 2568 954 2572
rect 1054 2568 1058 2572
rect 1174 2568 1178 2572
rect 1390 2568 1394 2572
rect 1518 2568 1522 2572
rect 2758 2568 2762 2572
rect 2782 2568 2786 2572
rect 2886 2568 2890 2572
rect 3174 2568 3178 2572
rect 3334 2568 3338 2572
rect 646 2558 650 2562
rect 654 2558 658 2562
rect 670 2558 674 2562
rect 718 2558 722 2562
rect 902 2558 906 2562
rect 910 2558 914 2562
rect 1278 2558 1282 2562
rect 1758 2558 1762 2562
rect 1774 2558 1778 2562
rect 1830 2558 1834 2562
rect 1910 2558 1914 2562
rect 2462 2558 2466 2562
rect 2502 2558 2506 2562
rect 2798 2558 2802 2562
rect 2838 2558 2842 2562
rect 2862 2558 2866 2562
rect 2870 2558 2874 2562
rect 3206 2558 3210 2562
rect 3230 2558 3234 2562
rect 158 2548 162 2552
rect 694 2548 698 2552
rect 806 2548 810 2552
rect 1382 2548 1386 2552
rect 1630 2548 1634 2552
rect 1806 2548 1810 2552
rect 1822 2548 1826 2552
rect 1934 2548 1938 2552
rect 2118 2548 2122 2552
rect 2502 2548 2506 2552
rect 2614 2548 2618 2552
rect 2734 2548 2738 2552
rect 2998 2548 3002 2552
rect 3174 2548 3178 2552
rect 3510 2548 3514 2552
rect 3614 2548 3618 2552
rect 3822 2548 3826 2552
rect 758 2538 762 2542
rect 878 2538 882 2542
rect 886 2538 890 2542
rect 974 2538 978 2542
rect 1102 2538 1106 2542
rect 1126 2538 1130 2542
rect 1142 2538 1146 2542
rect 1174 2538 1178 2542
rect 1478 2538 1482 2542
rect 1694 2538 1698 2542
rect 1734 2538 1738 2542
rect 1782 2538 1786 2542
rect 1846 2538 1850 2542
rect 2166 2538 2170 2542
rect 2462 2538 2466 2542
rect 2470 2538 2474 2542
rect 2894 2538 2898 2542
rect 3118 2538 3122 2542
rect 3126 2538 3130 2542
rect 3254 2538 3258 2542
rect 3734 2538 3738 2542
rect 382 2528 386 2532
rect 942 2528 946 2532
rect 1102 2528 1106 2532
rect 1222 2528 1226 2532
rect 1286 2528 1290 2532
rect 1622 2528 1626 2532
rect 1662 2528 1666 2532
rect 2150 2528 2154 2532
rect 2246 2528 2250 2532
rect 2598 2528 2602 2532
rect 2862 2528 2866 2532
rect 3214 2528 3218 2532
rect 3278 2528 3282 2532
rect 3382 2528 3386 2532
rect 3406 2528 3410 2532
rect 214 2518 218 2522
rect 782 2518 786 2522
rect 1206 2518 1210 2522
rect 1550 2518 1554 2522
rect 1822 2518 1826 2522
rect 1862 2518 1866 2522
rect 2078 2518 2082 2522
rect 2510 2518 2514 2522
rect 2606 2518 2610 2522
rect 2878 2518 2882 2522
rect 3494 2518 3498 2522
rect 3646 2518 3650 2522
rect 126 2508 130 2512
rect 462 2508 466 2512
rect 958 2508 962 2512
rect 982 2508 986 2512
rect 1190 2508 1194 2512
rect 1230 2508 1234 2512
rect 1542 2508 1546 2512
rect 1566 2508 1570 2512
rect 1782 2508 1786 2512
rect 2046 2508 2050 2512
rect 2406 2508 2410 2512
rect 2542 2508 2546 2512
rect 2678 2508 2682 2512
rect 2870 2508 2874 2512
rect 2878 2508 2882 2512
rect 3214 2508 3218 2512
rect 3222 2508 3226 2512
rect 3686 2508 3690 2512
rect 850 2503 854 2507
rect 858 2503 861 2507
rect 861 2503 862 2507
rect 1882 2503 1886 2507
rect 1890 2503 1893 2507
rect 1893 2503 1894 2507
rect 2906 2503 2910 2507
rect 2914 2503 2917 2507
rect 2917 2503 2918 2507
rect 934 2498 938 2502
rect 1462 2498 1466 2502
rect 1638 2498 1642 2502
rect 1670 2498 1674 2502
rect 2150 2498 2154 2502
rect 2422 2498 2426 2502
rect 2598 2498 2602 2502
rect 3022 2498 3026 2502
rect 1006 2488 1010 2492
rect 1206 2488 1210 2492
rect 1238 2488 1242 2492
rect 1510 2488 1514 2492
rect 1518 2488 1522 2492
rect 1918 2488 1922 2492
rect 2422 2488 2426 2492
rect 2582 2488 2586 2492
rect 2846 2488 2850 2492
rect 3222 2488 3226 2492
rect 3238 2488 3242 2492
rect 3270 2488 3274 2492
rect 3654 2488 3658 2492
rect 3678 2488 3682 2492
rect 238 2478 242 2482
rect 366 2478 370 2482
rect 638 2478 642 2482
rect 942 2478 946 2482
rect 982 2478 986 2482
rect 1830 2478 1834 2482
rect 2470 2478 2474 2482
rect 2606 2478 2610 2482
rect 2622 2478 2626 2482
rect 2822 2478 2826 2482
rect 2870 2478 2874 2482
rect 3134 2478 3138 2482
rect 3158 2478 3162 2482
rect 3246 2478 3250 2482
rect 3398 2478 3402 2482
rect 3566 2478 3570 2482
rect 3590 2478 3594 2482
rect 3742 2478 3746 2482
rect 190 2468 194 2472
rect 374 2468 378 2472
rect 534 2468 538 2472
rect 990 2468 994 2472
rect 1398 2468 1402 2472
rect 1470 2468 1474 2472
rect 1558 2468 1562 2472
rect 1958 2468 1962 2472
rect 2710 2468 2714 2472
rect 3062 2468 3066 2472
rect 3070 2468 3074 2472
rect 3150 2468 3154 2472
rect 3270 2468 3274 2472
rect 3390 2468 3394 2472
rect 3478 2468 3482 2472
rect 3750 2468 3754 2472
rect 62 2458 66 2462
rect 734 2458 738 2462
rect 830 2458 834 2462
rect 958 2458 962 2462
rect 1030 2458 1034 2462
rect 1070 2458 1074 2462
rect 1134 2458 1138 2462
rect 1198 2458 1202 2462
rect 1438 2458 1442 2462
rect 1510 2458 1514 2462
rect 1534 2458 1538 2462
rect 1942 2458 1946 2462
rect 1950 2458 1954 2462
rect 2654 2458 2658 2462
rect 2742 2458 2746 2462
rect 2854 2458 2858 2462
rect 2878 2458 2882 2462
rect 2950 2458 2954 2462
rect 3622 2458 3626 2462
rect 718 2448 722 2452
rect 934 2448 938 2452
rect 1838 2448 1842 2452
rect 1926 2448 1930 2452
rect 214 2438 218 2442
rect 2206 2448 2210 2452
rect 2462 2448 2466 2452
rect 2982 2448 2986 2452
rect 3350 2448 3354 2452
rect 3478 2448 3482 2452
rect 1134 2438 1138 2442
rect 1566 2438 1570 2442
rect 2310 2438 2314 2442
rect 2702 2438 2706 2442
rect 3022 2438 3026 2442
rect 3054 2438 3058 2442
rect 3438 2438 3442 2442
rect 3454 2438 3458 2442
rect 750 2428 754 2432
rect 1230 2428 1234 2432
rect 1542 2428 1546 2432
rect 1566 2428 1570 2432
rect 2302 2428 2306 2432
rect 2726 2428 2730 2432
rect 2782 2428 2786 2432
rect 206 2418 210 2422
rect 2102 2418 2106 2422
rect 3110 2418 3114 2422
rect 3622 2418 3626 2422
rect 1334 2408 1338 2412
rect 1814 2408 1818 2412
rect 2246 2408 2250 2412
rect 2590 2408 2594 2412
rect 3670 2408 3674 2412
rect 346 2403 350 2407
rect 354 2403 357 2407
rect 357 2403 358 2407
rect 1362 2403 1366 2407
rect 1370 2403 1373 2407
rect 1373 2403 1374 2407
rect 2386 2403 2390 2407
rect 2394 2403 2397 2407
rect 2397 2403 2398 2407
rect 3410 2403 3414 2407
rect 3418 2403 3421 2407
rect 3421 2403 3422 2407
rect 206 2398 210 2402
rect 966 2398 970 2402
rect 1470 2398 1474 2402
rect 1478 2398 1482 2402
rect 1774 2398 1778 2402
rect 2486 2398 2490 2402
rect 2990 2398 2994 2402
rect 3078 2398 3082 2402
rect 3382 2398 3386 2402
rect 790 2388 794 2392
rect 2422 2388 2426 2392
rect 2990 2388 2994 2392
rect 3462 2388 3466 2392
rect 494 2378 498 2382
rect 894 2378 898 2382
rect 1222 2378 1226 2382
rect 1590 2378 1594 2382
rect 3598 2378 3602 2382
rect 686 2368 690 2372
rect 1190 2368 1194 2372
rect 2614 2368 2618 2372
rect 3022 2368 3026 2372
rect 3198 2368 3202 2372
rect 3214 2368 3218 2372
rect 3478 2368 3482 2372
rect 3558 2368 3562 2372
rect 3742 2368 3746 2372
rect 742 2358 746 2362
rect 870 2358 874 2362
rect 1606 2358 1610 2362
rect 1670 2358 1674 2362
rect 1702 2358 1706 2362
rect 1782 2358 1786 2362
rect 2030 2358 2034 2362
rect 2358 2358 2362 2362
rect 2958 2358 2962 2362
rect 3446 2358 3450 2362
rect 3694 2358 3698 2362
rect 454 2348 458 2352
rect 646 2348 650 2352
rect 678 2348 682 2352
rect 894 2348 898 2352
rect 926 2348 930 2352
rect 990 2348 994 2352
rect 1118 2348 1122 2352
rect 1198 2348 1202 2352
rect 1382 2348 1386 2352
rect 1686 2348 1690 2352
rect 1838 2348 1842 2352
rect 1854 2348 1858 2352
rect 1958 2348 1962 2352
rect 2350 2348 2354 2352
rect 2838 2348 2842 2352
rect 2854 2348 2858 2352
rect 2894 2348 2898 2352
rect 3030 2348 3034 2352
rect 3134 2348 3138 2352
rect 3206 2348 3210 2352
rect 502 2338 506 2342
rect 1230 2338 1234 2342
rect 1294 2338 1298 2342
rect 1478 2338 1482 2342
rect 2310 2338 2314 2342
rect 2414 2338 2418 2342
rect 2742 2338 2746 2342
rect 2806 2338 2810 2342
rect 2846 2338 2850 2342
rect 2862 2338 2866 2342
rect 2870 2338 2874 2342
rect 2998 2338 3002 2342
rect 3062 2338 3066 2342
rect 3550 2338 3554 2342
rect 694 2328 698 2332
rect 1238 2328 1242 2332
rect 1262 2328 1266 2332
rect 1718 2328 1722 2332
rect 1814 2328 1818 2332
rect 2150 2328 2154 2332
rect 2342 2328 2346 2332
rect 2430 2328 2434 2332
rect 2438 2328 2442 2332
rect 2478 2328 2482 2332
rect 2790 2328 2794 2332
rect 2798 2328 2802 2332
rect 2830 2328 2834 2332
rect 3358 2328 3362 2332
rect 3494 2328 3498 2332
rect 870 2318 874 2322
rect 3094 2318 3098 2322
rect 3190 2318 3194 2322
rect 806 2308 810 2312
rect 838 2308 842 2312
rect 1846 2308 1850 2312
rect 1870 2308 1874 2312
rect 1942 2308 1946 2312
rect 2030 2308 2034 2312
rect 2926 2308 2930 2312
rect 3214 2308 3218 2312
rect 850 2303 854 2307
rect 858 2303 861 2307
rect 861 2303 862 2307
rect 1882 2303 1886 2307
rect 1890 2303 1893 2307
rect 1893 2303 1894 2307
rect 2906 2303 2910 2307
rect 2914 2303 2917 2307
rect 2917 2303 2918 2307
rect 462 2298 466 2302
rect 870 2298 874 2302
rect 2030 2298 2034 2302
rect 2846 2298 2850 2302
rect 3342 2298 3346 2302
rect 1854 2288 1858 2292
rect 2046 2288 2050 2292
rect 2422 2288 2426 2292
rect 3686 2288 3690 2292
rect 30 2278 34 2282
rect 1094 2278 1098 2282
rect 1110 2278 1114 2282
rect 1310 2278 1314 2282
rect 1734 2278 1738 2282
rect 1814 2278 1818 2282
rect 2118 2278 2122 2282
rect 2262 2278 2266 2282
rect 2470 2278 2474 2282
rect 2846 2278 2850 2282
rect 3118 2278 3122 2282
rect 3278 2278 3282 2282
rect 3438 2278 3442 2282
rect 3462 2278 3466 2282
rect 3542 2278 3546 2282
rect 3566 2278 3570 2282
rect 38 2268 42 2272
rect 1014 2268 1018 2272
rect 1446 2268 1450 2272
rect 1486 2268 1490 2272
rect 1502 2268 1506 2272
rect 1606 2268 1610 2272
rect 1790 2268 1794 2272
rect 1862 2268 1866 2272
rect 2006 2268 2010 2272
rect 2174 2268 2178 2272
rect 2374 2268 2378 2272
rect 2478 2268 2482 2272
rect 2630 2268 2634 2272
rect 2718 2268 2722 2272
rect 3038 2268 3042 2272
rect 3166 2268 3170 2272
rect 3206 2268 3210 2272
rect 3734 2268 3738 2272
rect 150 2258 154 2262
rect 198 2258 202 2262
rect 294 2258 298 2262
rect 822 2258 826 2262
rect 886 2258 890 2262
rect 1126 2258 1130 2262
rect 1294 2258 1298 2262
rect 1350 2258 1354 2262
rect 1382 2258 1386 2262
rect 1582 2258 1586 2262
rect 1750 2258 1754 2262
rect 2214 2258 2218 2262
rect 2294 2258 2298 2262
rect 2446 2258 2450 2262
rect 2542 2258 2546 2262
rect 2846 2258 2850 2262
rect 2982 2258 2986 2262
rect 3054 2258 3058 2262
rect 3198 2258 3202 2262
rect 3270 2258 3274 2262
rect 3318 2258 3322 2262
rect 3334 2258 3338 2262
rect 3694 2258 3698 2262
rect 3726 2258 3730 2262
rect 974 2248 978 2252
rect 1046 2248 1050 2252
rect 1062 2248 1066 2252
rect 1070 2248 1074 2252
rect 1510 2248 1514 2252
rect 1750 2248 1754 2252
rect 1846 2248 1850 2252
rect 2006 2248 2010 2252
rect 2086 2248 2090 2252
rect 2158 2248 2162 2252
rect 2614 2248 2618 2252
rect 3470 2248 3474 2252
rect 3566 2248 3570 2252
rect 614 2238 618 2242
rect 1038 2238 1042 2242
rect 1422 2238 1426 2242
rect 1526 2238 1530 2242
rect 1766 2238 1770 2242
rect 2278 2238 2282 2242
rect 2430 2238 2434 2242
rect 3038 2238 3042 2242
rect 3550 2238 3554 2242
rect 3662 2238 3666 2242
rect 1142 2228 1146 2232
rect 1206 2228 1210 2232
rect 2022 2228 2026 2232
rect 2174 2228 2178 2232
rect 286 2218 290 2222
rect 1814 2218 1818 2222
rect 1958 2218 1962 2222
rect 2006 2218 2010 2222
rect 2462 2218 2466 2222
rect 2822 2218 2826 2222
rect 2878 2218 2882 2222
rect 1166 2208 1170 2212
rect 1670 2208 1674 2212
rect 1734 2208 1738 2212
rect 1974 2208 1978 2212
rect 3222 2208 3226 2212
rect 346 2203 350 2207
rect 354 2203 357 2207
rect 357 2203 358 2207
rect 1362 2203 1366 2207
rect 1370 2203 1373 2207
rect 1373 2203 1374 2207
rect 2386 2203 2390 2207
rect 2394 2203 2397 2207
rect 2397 2203 2398 2207
rect 3410 2203 3414 2207
rect 3418 2203 3421 2207
rect 3421 2203 3422 2207
rect 2150 2198 2154 2202
rect 2222 2198 2226 2202
rect 2246 2198 2250 2202
rect 2606 2198 2610 2202
rect 3398 2198 3402 2202
rect 30 2188 34 2192
rect 422 2188 426 2192
rect 830 2188 834 2192
rect 1150 2188 1154 2192
rect 1518 2188 1522 2192
rect 2174 2188 2178 2192
rect 2598 2188 2602 2192
rect 2998 2188 3002 2192
rect 3030 2188 3034 2192
rect 3430 2188 3434 2192
rect 550 2178 554 2182
rect 574 2178 578 2182
rect 766 2178 770 2182
rect 1342 2178 1346 2182
rect 1502 2178 1506 2182
rect 1686 2178 1690 2182
rect 1718 2178 1722 2182
rect 1766 2178 1770 2182
rect 2662 2178 2666 2182
rect 3086 2178 3090 2182
rect 910 2168 914 2172
rect 1558 2168 1562 2172
rect 1814 2168 1818 2172
rect 1982 2168 1986 2172
rect 2022 2168 2026 2172
rect 2294 2168 2298 2172
rect 2462 2168 2466 2172
rect 2470 2168 2474 2172
rect 2510 2168 2514 2172
rect 3054 2168 3058 2172
rect 3606 2168 3610 2172
rect 734 2158 738 2162
rect 750 2158 754 2162
rect 798 2158 802 2162
rect 1102 2158 1106 2162
rect 1126 2158 1130 2162
rect 1854 2158 1858 2162
rect 1926 2158 1930 2162
rect 1966 2158 1970 2162
rect 2230 2158 2234 2162
rect 2430 2158 2434 2162
rect 2510 2158 2514 2162
rect 2526 2158 2530 2162
rect 2670 2158 2674 2162
rect 2686 2158 2690 2162
rect 3686 2158 3690 2162
rect 3694 2158 3698 2162
rect 526 2148 530 2152
rect 638 2148 642 2152
rect 710 2148 714 2152
rect 742 2148 746 2152
rect 1198 2148 1202 2152
rect 1270 2148 1274 2152
rect 1470 2148 1474 2152
rect 1550 2148 1554 2152
rect 1606 2148 1610 2152
rect 1614 2148 1618 2152
rect 2614 2148 2618 2152
rect 2654 2148 2658 2152
rect 2710 2148 2714 2152
rect 2782 2148 2786 2152
rect 2790 2148 2794 2152
rect 2814 2148 2818 2152
rect 2846 2148 2850 2152
rect 3598 2148 3602 2152
rect 3614 2148 3618 2152
rect 3710 2148 3714 2152
rect 134 2138 138 2142
rect 446 2138 450 2142
rect 526 2138 530 2142
rect 958 2138 962 2142
rect 1198 2138 1202 2142
rect 1310 2138 1314 2142
rect 1414 2138 1418 2142
rect 1910 2138 1914 2142
rect 2206 2138 2210 2142
rect 2446 2138 2450 2142
rect 2526 2138 2530 2142
rect 2718 2138 2722 2142
rect 2734 2138 2738 2142
rect 2750 2138 2754 2142
rect 2926 2138 2930 2142
rect 2958 2138 2962 2142
rect 3086 2138 3090 2142
rect 3158 2138 3162 2142
rect 3398 2138 3402 2142
rect 3622 2138 3626 2142
rect 366 2128 370 2132
rect 1254 2128 1258 2132
rect 1518 2128 1522 2132
rect 2094 2128 2098 2132
rect 2342 2128 2346 2132
rect 2438 2128 2442 2132
rect 2550 2128 2554 2132
rect 2606 2128 2610 2132
rect 2862 2128 2866 2132
rect 2878 2128 2882 2132
rect 2942 2128 2946 2132
rect 2958 2128 2962 2132
rect 3310 2128 3314 2132
rect 3326 2128 3330 2132
rect 3534 2128 3538 2132
rect 934 2118 938 2122
rect 1446 2118 1450 2122
rect 1454 2118 1458 2122
rect 1750 2118 1754 2122
rect 1870 2118 1874 2122
rect 1966 2118 1970 2122
rect 2214 2118 2218 2122
rect 2542 2118 2546 2122
rect 2590 2118 2594 2122
rect 2950 2118 2954 2122
rect 3110 2118 3114 2122
rect 3646 2118 3650 2122
rect 918 2108 922 2112
rect 1270 2108 1274 2112
rect 1310 2108 1314 2112
rect 1822 2108 1826 2112
rect 1862 2108 1866 2112
rect 2646 2108 2650 2112
rect 2894 2108 2898 2112
rect 3222 2108 3226 2112
rect 3238 2108 3242 2112
rect 3318 2108 3322 2112
rect 3350 2108 3354 2112
rect 850 2103 854 2107
rect 858 2103 861 2107
rect 861 2103 862 2107
rect 1882 2103 1886 2107
rect 1890 2103 1893 2107
rect 1893 2103 1894 2107
rect 2906 2103 2910 2107
rect 2914 2103 2917 2107
rect 2917 2103 2918 2107
rect 262 2098 266 2102
rect 718 2098 722 2102
rect 1614 2098 1618 2102
rect 1782 2098 1786 2102
rect 2206 2098 2210 2102
rect 2414 2098 2418 2102
rect 2494 2098 2498 2102
rect 2822 2098 2826 2102
rect 2926 2098 2930 2102
rect 3678 2098 3682 2102
rect 3774 2098 3778 2102
rect 1182 2088 1186 2092
rect 1590 2088 1594 2092
rect 1926 2088 1930 2092
rect 1958 2088 1962 2092
rect 1998 2088 2002 2092
rect 2430 2088 2434 2092
rect 2598 2088 2602 2092
rect 2622 2088 2626 2092
rect 2734 2088 2738 2092
rect 2806 2088 2810 2092
rect 2830 2088 2834 2092
rect 3750 2088 3754 2092
rect 1134 2078 1138 2082
rect 1278 2078 1282 2082
rect 1526 2078 1530 2082
rect 1622 2078 1626 2082
rect 1910 2078 1914 2082
rect 2182 2078 2186 2082
rect 2310 2078 2314 2082
rect 2422 2078 2426 2082
rect 2446 2078 2450 2082
rect 2782 2078 2786 2082
rect 2814 2078 2818 2082
rect 2830 2078 2834 2082
rect 3094 2078 3098 2082
rect 3374 2078 3378 2082
rect 3462 2078 3466 2082
rect 54 2068 58 2072
rect 230 2068 234 2072
rect 1878 2068 1882 2072
rect 2158 2068 2162 2072
rect 2566 2068 2570 2072
rect 2670 2068 2674 2072
rect 2926 2068 2930 2072
rect 3294 2068 3298 2072
rect 3302 2068 3306 2072
rect 3318 2068 3322 2072
rect 62 2058 66 2062
rect 1462 2058 1466 2062
rect 1582 2058 1586 2062
rect 1782 2058 1786 2062
rect 1798 2058 1802 2062
rect 1926 2058 1930 2062
rect 1974 2058 1978 2062
rect 2310 2058 2314 2062
rect 2470 2058 2474 2062
rect 2582 2058 2586 2062
rect 2614 2058 2618 2062
rect 2694 2058 2698 2062
rect 2774 2058 2778 2062
rect 3102 2058 3106 2062
rect 3126 2058 3130 2062
rect 3358 2058 3362 2062
rect 3446 2058 3450 2062
rect 3542 2058 3546 2062
rect 3622 2058 3626 2062
rect 470 2048 474 2052
rect 558 2048 562 2052
rect 630 2048 634 2052
rect 1390 2048 1394 2052
rect 1734 2048 1738 2052
rect 1798 2048 1802 2052
rect 1862 2048 1866 2052
rect 1942 2048 1946 2052
rect 2142 2048 2146 2052
rect 2182 2048 2186 2052
rect 2214 2048 2218 2052
rect 2350 2048 2354 2052
rect 2742 2048 2746 2052
rect 3046 2048 3050 2052
rect 3374 2048 3378 2052
rect 3566 2048 3570 2052
rect 3670 2048 3674 2052
rect 3734 2048 3738 2052
rect 454 2038 458 2042
rect 910 2038 914 2042
rect 1214 2038 1218 2042
rect 2006 2038 2010 2042
rect 2406 2038 2410 2042
rect 2438 2038 2442 2042
rect 2494 2038 2498 2042
rect 2598 2038 2602 2042
rect 2678 2038 2682 2042
rect 2894 2038 2898 2042
rect 2990 2038 2994 2042
rect 3126 2038 3130 2042
rect 3542 2038 3546 2042
rect 3646 2038 3650 2042
rect 3654 2038 3658 2042
rect 3734 2038 3738 2042
rect 230 2028 234 2032
rect 1774 2028 1778 2032
rect 2478 2028 2482 2032
rect 3366 2028 3370 2032
rect 3526 2028 3530 2032
rect 734 2018 738 2022
rect 1158 2018 1162 2022
rect 1566 2018 1570 2022
rect 1806 2018 1810 2022
rect 2934 2018 2938 2022
rect 3006 2018 3010 2022
rect 3294 2018 3298 2022
rect 3550 2018 3554 2022
rect 758 2008 762 2012
rect 950 2008 954 2012
rect 1174 2008 1178 2012
rect 1182 2008 1186 2012
rect 1838 2008 1842 2012
rect 2318 2008 2322 2012
rect 346 2003 350 2007
rect 354 2003 357 2007
rect 357 2003 358 2007
rect 1362 2003 1366 2007
rect 1370 2003 1373 2007
rect 1373 2003 1374 2007
rect 2386 2003 2390 2007
rect 2394 2003 2397 2007
rect 2397 2003 2398 2007
rect 3410 2003 3414 2007
rect 3418 2003 3421 2007
rect 3421 2003 3422 2007
rect 158 1998 162 2002
rect 1046 1998 1050 2002
rect 2230 1998 2234 2002
rect 2374 1998 2378 2002
rect 3398 1998 3402 2002
rect 886 1988 890 1992
rect 1030 1988 1034 1992
rect 1262 1988 1266 1992
rect 1318 1988 1322 1992
rect 1334 1988 1338 1992
rect 2150 1988 2154 1992
rect 2550 1988 2554 1992
rect 2838 1988 2842 1992
rect 2846 1988 2850 1992
rect 3142 1988 3146 1992
rect 3382 1988 3386 1992
rect 3390 1988 3394 1992
rect 526 1978 530 1982
rect 1198 1978 1202 1982
rect 566 1968 570 1972
rect 2366 1978 2370 1982
rect 2510 1978 2514 1982
rect 2518 1978 2522 1982
rect 2566 1978 2570 1982
rect 2774 1978 2778 1982
rect 1214 1968 1218 1972
rect 1294 1968 1298 1972
rect 2358 1968 2362 1972
rect 2462 1968 2466 1972
rect 2694 1968 2698 1972
rect 2870 1968 2874 1972
rect 3326 1968 3330 1972
rect 870 1958 874 1962
rect 998 1958 1002 1962
rect 1310 1958 1314 1962
rect 1710 1958 1714 1962
rect 1718 1958 1722 1962
rect 2206 1958 2210 1962
rect 2262 1958 2266 1962
rect 2454 1958 2458 1962
rect 2518 1958 2522 1962
rect 2574 1958 2578 1962
rect 3134 1958 3138 1962
rect 3390 1958 3394 1962
rect 3438 1958 3442 1962
rect 3590 1958 3594 1962
rect 3670 1958 3674 1962
rect 6 1948 10 1952
rect 62 1948 66 1952
rect 270 1948 274 1952
rect 638 1948 642 1952
rect 686 1948 690 1952
rect 726 1948 730 1952
rect 894 1948 898 1952
rect 990 1948 994 1952
rect 1382 1948 1386 1952
rect 1470 1948 1474 1952
rect 1534 1948 1538 1952
rect 1606 1948 1610 1952
rect 1686 1948 1690 1952
rect 1830 1948 1834 1952
rect 1846 1948 1850 1952
rect 1998 1948 2002 1952
rect 2406 1948 2410 1952
rect 2502 1948 2506 1952
rect 2614 1948 2618 1952
rect 2630 1948 2634 1952
rect 2710 1948 2714 1952
rect 2758 1948 2762 1952
rect 3022 1948 3026 1952
rect 3054 1948 3058 1952
rect 3062 1948 3066 1952
rect 3158 1948 3162 1952
rect 3302 1948 3306 1952
rect 46 1938 50 1942
rect 54 1938 58 1942
rect 190 1938 194 1942
rect 742 1938 746 1942
rect 918 1938 922 1942
rect 1622 1938 1626 1942
rect 1638 1938 1642 1942
rect 1974 1938 1978 1942
rect 2414 1938 2418 1942
rect 2430 1938 2434 1942
rect 2462 1938 2466 1942
rect 2566 1938 2570 1942
rect 2598 1938 2602 1942
rect 2622 1938 2626 1942
rect 2726 1938 2730 1942
rect 2974 1938 2978 1942
rect 3038 1938 3042 1942
rect 3150 1938 3154 1942
rect 3166 1938 3170 1942
rect 3286 1938 3290 1942
rect 3446 1938 3450 1942
rect 3758 1938 3762 1942
rect 478 1928 482 1932
rect 750 1928 754 1932
rect 1726 1928 1730 1932
rect 2030 1928 2034 1932
rect 2054 1928 2058 1932
rect 2126 1928 2130 1932
rect 2446 1928 2450 1932
rect 2478 1928 2482 1932
rect 2726 1928 2730 1932
rect 2750 1928 2754 1932
rect 2878 1928 2882 1932
rect 2966 1928 2970 1932
rect 3086 1928 3090 1932
rect 3094 1928 3098 1932
rect 3246 1928 3250 1932
rect 3510 1928 3514 1932
rect 3566 1928 3570 1932
rect 142 1918 146 1922
rect 494 1918 498 1922
rect 622 1918 626 1922
rect 774 1918 778 1922
rect 958 1918 962 1922
rect 1774 1918 1778 1922
rect 2710 1918 2714 1922
rect 2790 1918 2794 1922
rect 2894 1918 2898 1922
rect 2974 1918 2978 1922
rect 3446 1918 3450 1922
rect 110 1908 114 1912
rect 838 1908 842 1912
rect 950 1908 954 1912
rect 1582 1908 1586 1912
rect 1590 1908 1594 1912
rect 1950 1908 1954 1912
rect 1966 1908 1970 1912
rect 2118 1908 2122 1912
rect 2326 1908 2330 1912
rect 2406 1908 2410 1912
rect 2870 1908 2874 1912
rect 2934 1908 2938 1912
rect 2966 1908 2970 1912
rect 3166 1908 3170 1912
rect 3262 1908 3266 1912
rect 3414 1908 3418 1912
rect 850 1903 854 1907
rect 858 1903 861 1907
rect 861 1903 862 1907
rect 1882 1903 1886 1907
rect 1890 1903 1893 1907
rect 1893 1903 1894 1907
rect 790 1898 794 1902
rect 1526 1898 1530 1902
rect 1566 1898 1570 1902
rect 1806 1898 1810 1902
rect 2294 1898 2298 1902
rect 2906 1903 2910 1907
rect 2914 1903 2917 1907
rect 2917 1903 2918 1907
rect 2926 1898 2930 1902
rect 3038 1898 3042 1902
rect 3054 1898 3058 1902
rect 3086 1898 3090 1902
rect 3222 1898 3226 1902
rect 3278 1898 3282 1902
rect 3310 1898 3314 1902
rect 958 1888 962 1892
rect 1590 1888 1594 1892
rect 1598 1888 1602 1892
rect 1702 1888 1706 1892
rect 1742 1888 1746 1892
rect 2286 1888 2290 1892
rect 2430 1888 2434 1892
rect 2686 1888 2690 1892
rect 2774 1888 2778 1892
rect 3342 1888 3346 1892
rect 3566 1888 3570 1892
rect 3654 1888 3658 1892
rect 126 1878 130 1882
rect 550 1878 554 1882
rect 694 1878 698 1882
rect 702 1878 706 1882
rect 1062 1878 1066 1882
rect 1198 1878 1202 1882
rect 1302 1878 1306 1882
rect 1662 1878 1666 1882
rect 1726 1878 1730 1882
rect 2102 1878 2106 1882
rect 2270 1878 2274 1882
rect 2438 1878 2442 1882
rect 2662 1878 2666 1882
rect 2838 1878 2842 1882
rect 2918 1878 2922 1882
rect 3382 1878 3386 1882
rect 3478 1878 3482 1882
rect 270 1868 274 1872
rect 510 1868 514 1872
rect 918 1868 922 1872
rect 966 1868 970 1872
rect 1190 1868 1194 1872
rect 1334 1868 1338 1872
rect 1510 1868 1514 1872
rect 1518 1868 1522 1872
rect 2174 1868 2178 1872
rect 2198 1868 2202 1872
rect 2302 1868 2306 1872
rect 2366 1868 2370 1872
rect 3190 1868 3194 1872
rect 3758 1868 3762 1872
rect 454 1858 458 1862
rect 590 1858 594 1862
rect 630 1858 634 1862
rect 726 1858 730 1862
rect 782 1858 786 1862
rect 1070 1858 1074 1862
rect 1238 1858 1242 1862
rect 1302 1858 1306 1862
rect 1430 1858 1434 1862
rect 2342 1858 2346 1862
rect 2414 1858 2418 1862
rect 2454 1858 2458 1862
rect 2526 1858 2530 1862
rect 2558 1858 2562 1862
rect 2766 1858 2770 1862
rect 2870 1858 2874 1862
rect 2942 1858 2946 1862
rect 2982 1858 2986 1862
rect 3118 1858 3122 1862
rect 3262 1858 3266 1862
rect 3342 1858 3346 1862
rect 3374 1858 3378 1862
rect 6 1848 10 1852
rect 614 1848 618 1852
rect 774 1848 778 1852
rect 1686 1848 1690 1852
rect 2350 1848 2354 1852
rect 2646 1848 2650 1852
rect 2766 1848 2770 1852
rect 3302 1848 3306 1852
rect 3526 1848 3530 1852
rect 3558 1848 3562 1852
rect 3590 1848 3594 1852
rect 3750 1848 3754 1852
rect 566 1838 570 1842
rect 942 1838 946 1842
rect 1182 1838 1186 1842
rect 1654 1838 1658 1842
rect 1950 1838 1954 1842
rect 2262 1838 2266 1842
rect 2406 1838 2410 1842
rect 2454 1838 2458 1842
rect 3254 1838 3258 1842
rect 3390 1838 3394 1842
rect 3694 1838 3698 1842
rect 3734 1838 3738 1842
rect 654 1828 658 1832
rect 1150 1828 1154 1832
rect 1582 1828 1586 1832
rect 2566 1828 2570 1832
rect 3102 1828 3106 1832
rect 3150 1828 3154 1832
rect 3758 1828 3762 1832
rect 806 1818 810 1822
rect 1574 1818 1578 1822
rect 2358 1818 2362 1822
rect 2854 1818 2858 1822
rect 3270 1818 3274 1822
rect 3390 1818 3394 1822
rect 1182 1808 1186 1812
rect 1550 1808 1554 1812
rect 2406 1808 2410 1812
rect 3022 1808 3026 1812
rect 3062 1808 3066 1812
rect 346 1803 350 1807
rect 354 1803 357 1807
rect 357 1803 358 1807
rect 1362 1803 1366 1807
rect 1370 1803 1373 1807
rect 1373 1803 1374 1807
rect 2386 1803 2390 1807
rect 2394 1803 2397 1807
rect 2397 1803 2398 1807
rect 3410 1803 3414 1807
rect 3418 1803 3421 1807
rect 3421 1803 3422 1807
rect 878 1798 882 1802
rect 1086 1798 1090 1802
rect 1574 1798 1578 1802
rect 2782 1798 2786 1802
rect 3542 1798 3546 1802
rect 3590 1798 3594 1802
rect 750 1788 754 1792
rect 1278 1788 1282 1792
rect 2334 1788 2338 1792
rect 2430 1788 2434 1792
rect 3238 1788 3242 1792
rect 3598 1788 3602 1792
rect 718 1778 722 1782
rect 1590 1778 1594 1782
rect 1670 1778 1674 1782
rect 1766 1778 1770 1782
rect 1798 1778 1802 1782
rect 2278 1778 2282 1782
rect 2318 1778 2322 1782
rect 1910 1768 1914 1772
rect 2118 1768 2122 1772
rect 2462 1768 2466 1772
rect 2510 1768 2514 1772
rect 2574 1768 2578 1772
rect 2710 1768 2714 1772
rect 2758 1768 2762 1772
rect 2950 1768 2954 1772
rect 3222 1768 3226 1772
rect 3382 1768 3386 1772
rect 798 1758 802 1762
rect 958 1758 962 1762
rect 1790 1758 1794 1762
rect 1806 1758 1810 1762
rect 2070 1758 2074 1762
rect 2382 1758 2386 1762
rect 2526 1758 2530 1762
rect 2870 1758 2874 1762
rect 3190 1758 3194 1762
rect 3286 1758 3290 1762
rect 3534 1758 3538 1762
rect 3646 1758 3650 1762
rect 294 1748 298 1752
rect 310 1748 314 1752
rect 382 1748 386 1752
rect 478 1748 482 1752
rect 534 1748 538 1752
rect 670 1748 674 1752
rect 790 1748 794 1752
rect 814 1748 818 1752
rect 1382 1748 1386 1752
rect 1606 1748 1610 1752
rect 2630 1748 2634 1752
rect 2670 1748 2674 1752
rect 2758 1748 2762 1752
rect 2862 1748 2866 1752
rect 2870 1748 2874 1752
rect 3070 1748 3074 1752
rect 3166 1748 3170 1752
rect 3430 1748 3434 1752
rect 3462 1748 3466 1752
rect 3518 1748 3522 1752
rect 3670 1748 3674 1752
rect 3750 1748 3754 1752
rect 134 1738 138 1742
rect 462 1738 466 1742
rect 662 1738 666 1742
rect 806 1738 810 1742
rect 1046 1738 1050 1742
rect 1222 1738 1226 1742
rect 1374 1738 1378 1742
rect 1574 1738 1578 1742
rect 1582 1738 1586 1742
rect 1646 1738 1650 1742
rect 1654 1738 1658 1742
rect 1982 1738 1986 1742
rect 2294 1738 2298 1742
rect 2366 1738 2370 1742
rect 2374 1738 2378 1742
rect 2526 1738 2530 1742
rect 2566 1738 2570 1742
rect 2686 1738 2690 1742
rect 2702 1738 2706 1742
rect 2718 1738 2722 1742
rect 2814 1738 2818 1742
rect 3126 1738 3130 1742
rect 3702 1738 3706 1742
rect 126 1728 130 1732
rect 294 1728 298 1732
rect 374 1728 378 1732
rect 414 1728 418 1732
rect 422 1728 426 1732
rect 438 1728 442 1732
rect 686 1728 690 1732
rect 774 1728 778 1732
rect 950 1728 954 1732
rect 1030 1728 1034 1732
rect 1062 1728 1066 1732
rect 1622 1728 1626 1732
rect 1694 1728 1698 1732
rect 1902 1728 1906 1732
rect 1990 1728 1994 1732
rect 2486 1728 2490 1732
rect 2550 1728 2554 1732
rect 2646 1728 2650 1732
rect 2718 1728 2722 1732
rect 2990 1728 2994 1732
rect 3278 1728 3282 1732
rect 3438 1728 3442 1732
rect 3694 1728 3698 1732
rect 542 1718 546 1722
rect 934 1718 938 1722
rect 1022 1718 1026 1722
rect 1038 1718 1042 1722
rect 1918 1718 1922 1722
rect 2126 1718 2130 1722
rect 2958 1718 2962 1722
rect 2966 1718 2970 1722
rect 3054 1718 3058 1722
rect 3646 1718 3650 1722
rect 366 1708 370 1712
rect 782 1708 786 1712
rect 878 1708 882 1712
rect 966 1708 970 1712
rect 1638 1708 1642 1712
rect 1910 1708 1914 1712
rect 2398 1708 2402 1712
rect 2886 1708 2890 1712
rect 2990 1708 2994 1712
rect 3078 1708 3082 1712
rect 3102 1708 3106 1712
rect 3542 1708 3546 1712
rect 3646 1708 3650 1712
rect 850 1703 854 1707
rect 858 1703 861 1707
rect 861 1703 862 1707
rect 1882 1703 1886 1707
rect 1890 1703 1893 1707
rect 1893 1703 1894 1707
rect 2906 1703 2910 1707
rect 2914 1703 2917 1707
rect 2917 1703 2918 1707
rect 462 1698 466 1702
rect 502 1698 506 1702
rect 1870 1698 1874 1702
rect 1902 1698 1906 1702
rect 2134 1698 2138 1702
rect 2958 1698 2962 1702
rect 3230 1698 3234 1702
rect 390 1688 394 1692
rect 902 1688 906 1692
rect 1062 1688 1066 1692
rect 1230 1688 1234 1692
rect 1478 1688 1482 1692
rect 1774 1688 1778 1692
rect 1910 1688 1914 1692
rect 2062 1688 2066 1692
rect 2374 1688 2378 1692
rect 2550 1688 2554 1692
rect 2710 1688 2714 1692
rect 2718 1688 2722 1692
rect 94 1678 98 1682
rect 502 1678 506 1682
rect 662 1678 666 1682
rect 1238 1678 1242 1682
rect 1518 1678 1522 1682
rect 1638 1678 1642 1682
rect 2230 1678 2234 1682
rect 2294 1678 2298 1682
rect 2486 1678 2490 1682
rect 2998 1688 3002 1692
rect 2742 1678 2746 1682
rect 2846 1678 2850 1682
rect 3006 1678 3010 1682
rect 3070 1678 3074 1682
rect 3310 1678 3314 1682
rect 3398 1678 3402 1682
rect 3526 1678 3530 1682
rect 6 1668 10 1672
rect 110 1668 114 1672
rect 238 1668 242 1672
rect 334 1668 338 1672
rect 718 1668 722 1672
rect 830 1668 834 1672
rect 1014 1668 1018 1672
rect 1038 1668 1042 1672
rect 1110 1668 1114 1672
rect 1182 1668 1186 1672
rect 1238 1668 1242 1672
rect 1486 1668 1490 1672
rect 1510 1668 1514 1672
rect 1590 1668 1594 1672
rect 1726 1668 1730 1672
rect 1782 1668 1786 1672
rect 1918 1668 1922 1672
rect 2094 1668 2098 1672
rect 2406 1668 2410 1672
rect 2846 1668 2850 1672
rect 3174 1668 3178 1672
rect 3230 1668 3234 1672
rect 3318 1668 3322 1672
rect 3518 1668 3522 1672
rect 3750 1668 3754 1672
rect 750 1658 754 1662
rect 798 1658 802 1662
rect 886 1658 890 1662
rect 942 1658 946 1662
rect 982 1658 986 1662
rect 990 1658 994 1662
rect 1102 1658 1106 1662
rect 1342 1658 1346 1662
rect 1350 1658 1354 1662
rect 1382 1658 1386 1662
rect 1670 1658 1674 1662
rect 1774 1658 1778 1662
rect 1806 1658 1810 1662
rect 2486 1658 2490 1662
rect 2686 1658 2690 1662
rect 2774 1658 2778 1662
rect 2822 1658 2826 1662
rect 3134 1658 3138 1662
rect 3694 1658 3698 1662
rect 3734 1658 3738 1662
rect 678 1648 682 1652
rect 870 1648 874 1652
rect 998 1648 1002 1652
rect 1454 1648 1458 1652
rect 1750 1648 1754 1652
rect 2350 1648 2354 1652
rect 2374 1648 2378 1652
rect 2574 1648 2578 1652
rect 3158 1648 3162 1652
rect 3750 1648 3754 1652
rect 526 1638 530 1642
rect 1334 1638 1338 1642
rect 1782 1638 1786 1642
rect 2686 1638 2690 1642
rect 3046 1638 3050 1642
rect 3238 1638 3242 1642
rect 3574 1638 3578 1642
rect 3670 1638 3674 1642
rect 518 1628 522 1632
rect 838 1628 842 1632
rect 1182 1628 1186 1632
rect 534 1618 538 1622
rect 1302 1618 1306 1622
rect 1326 1618 1330 1622
rect 3302 1618 3306 1622
rect 3558 1618 3562 1622
rect 750 1608 754 1612
rect 766 1608 770 1612
rect 918 1608 922 1612
rect 1254 1608 1258 1612
rect 1646 1608 1650 1612
rect 1654 1608 1658 1612
rect 1846 1608 1850 1612
rect 1926 1608 1930 1612
rect 3078 1608 3082 1612
rect 3086 1608 3090 1612
rect 346 1603 350 1607
rect 354 1603 357 1607
rect 357 1603 358 1607
rect 1362 1603 1366 1607
rect 1370 1603 1373 1607
rect 1373 1603 1374 1607
rect 2386 1603 2390 1607
rect 2394 1603 2397 1607
rect 2397 1603 2398 1607
rect 3410 1603 3414 1607
rect 3418 1603 3421 1607
rect 3421 1603 3422 1607
rect 1030 1598 1034 1602
rect 1238 1598 1242 1602
rect 1350 1598 1354 1602
rect 1614 1598 1618 1602
rect 1662 1598 1666 1602
rect 2366 1598 2370 1602
rect 2830 1598 2834 1602
rect 3486 1598 3490 1602
rect 3646 1598 3650 1602
rect 726 1588 730 1592
rect 1286 1588 1290 1592
rect 1630 1588 1634 1592
rect 2038 1588 2042 1592
rect 3734 1588 3738 1592
rect 1150 1578 1154 1582
rect 1446 1578 1450 1582
rect 1486 1578 1490 1582
rect 1862 1578 1866 1582
rect 2662 1578 2666 1582
rect 3142 1578 3146 1582
rect 3446 1578 3450 1582
rect 3486 1578 3490 1582
rect 742 1568 746 1572
rect 2230 1568 2234 1572
rect 3046 1568 3050 1572
rect 3222 1568 3226 1572
rect 3510 1568 3514 1572
rect 3758 1568 3762 1572
rect 302 1558 306 1562
rect 470 1558 474 1562
rect 1086 1558 1090 1562
rect 1902 1558 1906 1562
rect 2054 1558 2058 1562
rect 2734 1558 2738 1562
rect 2798 1558 2802 1562
rect 3086 1558 3090 1562
rect 3126 1558 3130 1562
rect 3246 1558 3250 1562
rect 3286 1558 3290 1562
rect 6 1548 10 1552
rect 822 1548 826 1552
rect 926 1548 930 1552
rect 1614 1548 1618 1552
rect 1742 1548 1746 1552
rect 2526 1548 2530 1552
rect 2598 1548 2602 1552
rect 3270 1548 3274 1552
rect 3350 1548 3354 1552
rect 3478 1548 3482 1552
rect 3510 1548 3514 1552
rect 3654 1548 3658 1552
rect 3710 1548 3714 1552
rect 3726 1548 3730 1552
rect 462 1538 466 1542
rect 670 1538 674 1542
rect 1790 1538 1794 1542
rect 1798 1538 1802 1542
rect 2126 1538 2130 1542
rect 2830 1538 2834 1542
rect 3230 1538 3234 1542
rect 3310 1538 3314 1542
rect 3382 1538 3386 1542
rect 462 1528 466 1532
rect 806 1528 810 1532
rect 950 1528 954 1532
rect 1190 1528 1194 1532
rect 1206 1528 1210 1532
rect 1870 1528 1874 1532
rect 2022 1528 2026 1532
rect 2502 1528 2506 1532
rect 3238 1528 3242 1532
rect 3262 1528 3266 1532
rect 3550 1528 3554 1532
rect 6 1518 10 1522
rect 1326 1518 1330 1522
rect 1446 1518 1450 1522
rect 1718 1518 1722 1522
rect 2870 1518 2874 1522
rect 3062 1518 3066 1522
rect 3238 1518 3242 1522
rect 430 1508 434 1512
rect 718 1508 722 1512
rect 830 1508 834 1512
rect 942 1508 946 1512
rect 1174 1508 1178 1512
rect 1278 1508 1282 1512
rect 1742 1508 1746 1512
rect 2710 1508 2714 1512
rect 2814 1508 2818 1512
rect 3070 1508 3074 1512
rect 3302 1508 3306 1512
rect 3310 1508 3314 1512
rect 3334 1508 3338 1512
rect 3350 1508 3354 1512
rect 850 1503 854 1507
rect 858 1503 861 1507
rect 861 1503 862 1507
rect 1882 1503 1886 1507
rect 1890 1503 1893 1507
rect 1893 1503 1894 1507
rect 2906 1503 2910 1507
rect 2914 1503 2917 1507
rect 2917 1503 2918 1507
rect 646 1498 650 1502
rect 1454 1498 1458 1502
rect 2862 1498 2866 1502
rect 3110 1498 3114 1502
rect 734 1488 738 1492
rect 846 1488 850 1492
rect 990 1488 994 1492
rect 1094 1488 1098 1492
rect 1110 1488 1114 1492
rect 1166 1488 1170 1492
rect 1182 1488 1186 1492
rect 1350 1488 1354 1492
rect 1950 1488 1954 1492
rect 1966 1488 1970 1492
rect 2174 1488 2178 1492
rect 2598 1488 2602 1492
rect 2718 1488 2722 1492
rect 3022 1488 3026 1492
rect 3214 1488 3218 1492
rect 3614 1488 3618 1492
rect 238 1478 242 1482
rect 390 1478 394 1482
rect 518 1478 522 1482
rect 654 1478 658 1482
rect 1310 1478 1314 1482
rect 1902 1478 1906 1482
rect 1910 1478 1914 1482
rect 2574 1478 2578 1482
rect 2758 1478 2762 1482
rect 2838 1478 2842 1482
rect 3158 1478 3162 1482
rect 3262 1478 3266 1482
rect 3542 1478 3546 1482
rect 3574 1478 3578 1482
rect 3694 1478 3698 1482
rect 422 1468 426 1472
rect 838 1468 842 1472
rect 1054 1468 1058 1472
rect 2590 1468 2594 1472
rect 2598 1468 2602 1472
rect 798 1458 802 1462
rect 966 1458 970 1462
rect 1062 1458 1066 1462
rect 1134 1458 1138 1462
rect 1206 1458 1210 1462
rect 1318 1458 1322 1462
rect 1558 1458 1562 1462
rect 1798 1458 1802 1462
rect 1910 1458 1914 1462
rect 2038 1458 2042 1462
rect 2414 1458 2418 1462
rect 2502 1458 2506 1462
rect 2678 1468 2682 1472
rect 2846 1468 2850 1472
rect 3014 1468 3018 1472
rect 3174 1468 3178 1472
rect 3462 1468 3466 1472
rect 3486 1468 3490 1472
rect 3694 1468 3698 1472
rect 2726 1458 2730 1462
rect 2998 1458 3002 1462
rect 3158 1458 3162 1462
rect 3454 1458 3458 1462
rect 3462 1458 3466 1462
rect 3534 1458 3538 1462
rect 3598 1458 3602 1462
rect 3774 1458 3778 1462
rect 494 1448 498 1452
rect 590 1448 594 1452
rect 1014 1448 1018 1452
rect 1446 1448 1450 1452
rect 1550 1448 1554 1452
rect 1630 1448 1634 1452
rect 1878 1448 1882 1452
rect 1942 1448 1946 1452
rect 2062 1448 2066 1452
rect 2310 1448 2314 1452
rect 2366 1448 2370 1452
rect 2470 1448 2474 1452
rect 2806 1448 2810 1452
rect 2950 1448 2954 1452
rect 3150 1448 3154 1452
rect 3374 1448 3378 1452
rect 3622 1448 3626 1452
rect 3694 1448 3698 1452
rect 3774 1448 3778 1452
rect 1278 1438 1282 1442
rect 2078 1438 2082 1442
rect 2422 1438 2426 1442
rect 2694 1438 2698 1442
rect 782 1428 786 1432
rect 2798 1428 2802 1432
rect 3646 1428 3650 1432
rect 166 1418 170 1422
rect 182 1418 186 1422
rect 750 1418 754 1422
rect 1078 1418 1082 1422
rect 1382 1418 1386 1422
rect 2422 1418 2426 1422
rect 3054 1418 3058 1422
rect 3126 1418 3130 1422
rect 2694 1408 2698 1412
rect 2798 1408 2802 1412
rect 3006 1408 3010 1412
rect 3014 1408 3018 1412
rect 3630 1408 3634 1412
rect 346 1403 350 1407
rect 354 1403 357 1407
rect 357 1403 358 1407
rect 1362 1403 1366 1407
rect 1370 1403 1373 1407
rect 1373 1403 1374 1407
rect 2386 1403 2390 1407
rect 2394 1403 2397 1407
rect 2397 1403 2398 1407
rect 566 1398 570 1402
rect 582 1398 586 1402
rect 934 1398 938 1402
rect 1350 1398 1354 1402
rect 1622 1398 1626 1402
rect 1790 1398 1794 1402
rect 2222 1398 2226 1402
rect 3410 1403 3414 1407
rect 3418 1403 3421 1407
rect 3421 1403 3422 1407
rect 3110 1398 3114 1402
rect 3150 1398 3154 1402
rect 3286 1398 3290 1402
rect 3582 1398 3586 1402
rect 510 1388 514 1392
rect 670 1388 674 1392
rect 758 1388 762 1392
rect 806 1388 810 1392
rect 1494 1388 1498 1392
rect 1886 1388 1890 1392
rect 3486 1388 3490 1392
rect 3726 1388 3730 1392
rect 886 1378 890 1382
rect 1038 1378 1042 1382
rect 1174 1378 1178 1382
rect 1606 1378 1610 1382
rect 2846 1378 2850 1382
rect 2886 1378 2890 1382
rect 3014 1378 3018 1382
rect 3134 1378 3138 1382
rect 3326 1378 3330 1382
rect 382 1368 386 1372
rect 2270 1368 2274 1372
rect 2510 1368 2514 1372
rect 2958 1368 2962 1372
rect 3110 1368 3114 1372
rect 3246 1368 3250 1372
rect 3630 1368 3634 1372
rect 182 1358 186 1362
rect 838 1358 842 1362
rect 942 1358 946 1362
rect 1126 1358 1130 1362
rect 1454 1358 1458 1362
rect 1678 1358 1682 1362
rect 1774 1358 1778 1362
rect 1878 1358 1882 1362
rect 2078 1358 2082 1362
rect 2166 1358 2170 1362
rect 2326 1358 2330 1362
rect 2502 1358 2506 1362
rect 2790 1358 2794 1362
rect 2878 1358 2882 1362
rect 3342 1358 3346 1362
rect 3510 1358 3514 1362
rect 3614 1358 3618 1362
rect 3670 1358 3674 1362
rect 3774 1358 3778 1362
rect 302 1348 306 1352
rect 470 1348 474 1352
rect 846 1348 850 1352
rect 1270 1348 1274 1352
rect 1430 1348 1434 1352
rect 1470 1348 1474 1352
rect 2094 1348 2098 1352
rect 2190 1348 2194 1352
rect 2262 1348 2266 1352
rect 3206 1348 3210 1352
rect 3334 1348 3338 1352
rect 3526 1348 3530 1352
rect 3542 1348 3546 1352
rect 3598 1348 3602 1352
rect 3646 1348 3650 1352
rect 6 1338 10 1342
rect 174 1338 178 1342
rect 566 1338 570 1342
rect 886 1338 890 1342
rect 950 1338 954 1342
rect 1070 1338 1074 1342
rect 1262 1338 1266 1342
rect 1310 1338 1314 1342
rect 2278 1338 2282 1342
rect 2374 1338 2378 1342
rect 2790 1338 2794 1342
rect 2862 1338 2866 1342
rect 3318 1338 3322 1342
rect 3374 1338 3378 1342
rect 3446 1338 3450 1342
rect 542 1328 546 1332
rect 574 1328 578 1332
rect 830 1328 834 1332
rect 1014 1328 1018 1332
rect 1246 1328 1250 1332
rect 1406 1328 1410 1332
rect 1614 1328 1618 1332
rect 1702 1328 1706 1332
rect 1718 1328 1722 1332
rect 2062 1328 2066 1332
rect 2134 1328 2138 1332
rect 2150 1328 2154 1332
rect 2238 1328 2242 1332
rect 2454 1328 2458 1332
rect 2678 1328 2682 1332
rect 2870 1328 2874 1332
rect 2966 1328 2970 1332
rect 3110 1328 3114 1332
rect 3222 1328 3226 1332
rect 3614 1328 3618 1332
rect 3646 1328 3650 1332
rect 478 1318 482 1322
rect 486 1318 490 1322
rect 694 1318 698 1322
rect 1910 1318 1914 1322
rect 2526 1318 2530 1322
rect 3094 1318 3098 1322
rect 3134 1318 3138 1322
rect 3158 1318 3162 1322
rect 3358 1318 3362 1322
rect 3462 1318 3466 1322
rect 3502 1318 3506 1322
rect 3686 1318 3690 1322
rect 526 1308 530 1312
rect 886 1308 890 1312
rect 1062 1308 1066 1312
rect 1094 1308 1098 1312
rect 1558 1308 1562 1312
rect 1934 1308 1938 1312
rect 2926 1308 2930 1312
rect 3086 1308 3090 1312
rect 850 1303 854 1307
rect 858 1303 861 1307
rect 861 1303 862 1307
rect 1882 1303 1886 1307
rect 1890 1303 1893 1307
rect 1893 1303 1894 1307
rect 2906 1303 2910 1307
rect 2914 1303 2917 1307
rect 2917 1303 2918 1307
rect 670 1298 674 1302
rect 894 1298 898 1302
rect 1094 1298 1098 1302
rect 1142 1298 1146 1302
rect 1830 1298 1834 1302
rect 2342 1298 2346 1302
rect 3174 1298 3178 1302
rect 438 1288 442 1292
rect 462 1288 466 1292
rect 734 1288 738 1292
rect 2086 1288 2090 1292
rect 2126 1288 2130 1292
rect 2270 1288 2274 1292
rect 2582 1288 2586 1292
rect 2822 1288 2826 1292
rect 2990 1288 2994 1292
rect 3286 1288 3290 1292
rect 3358 1288 3362 1292
rect 3686 1288 3690 1292
rect 382 1278 386 1282
rect 958 1278 962 1282
rect 1902 1278 1906 1282
rect 38 1268 42 1272
rect 486 1268 490 1272
rect 2294 1278 2298 1282
rect 2350 1278 2354 1282
rect 2446 1278 2450 1282
rect 2630 1278 2634 1282
rect 2678 1278 2682 1282
rect 3062 1278 3066 1282
rect 3134 1278 3138 1282
rect 3214 1278 3218 1282
rect 3310 1278 3314 1282
rect 1110 1268 1114 1272
rect 1134 1268 1138 1272
rect 1150 1268 1154 1272
rect 1286 1268 1290 1272
rect 1662 1268 1666 1272
rect 1694 1268 1698 1272
rect 1726 1268 1730 1272
rect 1846 1268 1850 1272
rect 1942 1268 1946 1272
rect 2238 1268 2242 1272
rect 2374 1268 2378 1272
rect 2782 1268 2786 1272
rect 3006 1268 3010 1272
rect 3342 1268 3346 1272
rect 3422 1268 3426 1272
rect 3486 1268 3490 1272
rect 3510 1268 3514 1272
rect 1078 1258 1082 1262
rect 1718 1258 1722 1262
rect 2246 1258 2250 1262
rect 2518 1258 2522 1262
rect 2542 1258 2546 1262
rect 2566 1258 2570 1262
rect 2614 1258 2618 1262
rect 2654 1258 2658 1262
rect 2758 1258 2762 1262
rect 2950 1258 2954 1262
rect 2966 1258 2970 1262
rect 3086 1258 3090 1262
rect 3166 1258 3170 1262
rect 3558 1258 3562 1262
rect 3630 1258 3634 1262
rect 3686 1258 3690 1262
rect 3750 1258 3754 1262
rect 774 1248 778 1252
rect 1198 1248 1202 1252
rect 1278 1248 1282 1252
rect 1646 1248 1650 1252
rect 2534 1248 2538 1252
rect 2982 1248 2986 1252
rect 3078 1248 3082 1252
rect 3230 1248 3234 1252
rect 3574 1248 3578 1252
rect 3582 1248 3586 1252
rect 3598 1248 3602 1252
rect 166 1238 170 1242
rect 262 1238 266 1242
rect 1998 1238 2002 1242
rect 2622 1238 2626 1242
rect 3238 1238 3242 1242
rect 3622 1238 3626 1242
rect 3670 1238 3674 1242
rect 3686 1238 3690 1242
rect 3750 1238 3754 1242
rect 622 1228 626 1232
rect 1118 1228 1122 1232
rect 2990 1228 2994 1232
rect 1462 1218 1466 1222
rect 1742 1218 1746 1222
rect 2038 1218 2042 1222
rect 2222 1218 2226 1222
rect 2318 1218 2322 1222
rect 1118 1208 1122 1212
rect 2406 1208 2410 1212
rect 2526 1208 2530 1212
rect 3182 1208 3186 1212
rect 3478 1208 3482 1212
rect 346 1203 350 1207
rect 354 1203 357 1207
rect 357 1203 358 1207
rect 638 1198 642 1202
rect 1362 1203 1366 1207
rect 1370 1203 1373 1207
rect 1373 1203 1374 1207
rect 2386 1203 2390 1207
rect 2394 1203 2397 1207
rect 2397 1203 2398 1207
rect 3410 1203 3414 1207
rect 3418 1203 3421 1207
rect 3421 1203 3422 1207
rect 1134 1198 1138 1202
rect 1382 1198 1386 1202
rect 1766 1198 1770 1202
rect 2638 1198 2642 1202
rect 3230 1198 3234 1202
rect 1270 1188 1274 1192
rect 1926 1188 1930 1192
rect 1974 1188 1978 1192
rect 2742 1188 2746 1192
rect 3358 1188 3362 1192
rect 3758 1188 3762 1192
rect 430 1178 434 1182
rect 686 1178 690 1182
rect 886 1178 890 1182
rect 1350 1178 1354 1182
rect 1726 1178 1730 1182
rect 1774 1178 1778 1182
rect 1806 1178 1810 1182
rect 1814 1178 1818 1182
rect 2334 1178 2338 1182
rect 2462 1178 2466 1182
rect 2942 1178 2946 1182
rect 6 1168 10 1172
rect 230 1168 234 1172
rect 454 1168 458 1172
rect 510 1168 514 1172
rect 566 1168 570 1172
rect 1326 1168 1330 1172
rect 2302 1168 2306 1172
rect 2422 1168 2426 1172
rect 2486 1168 2490 1172
rect 2606 1168 2610 1172
rect 2782 1168 2786 1172
rect 2806 1168 2810 1172
rect 2942 1168 2946 1172
rect 3542 1168 3546 1172
rect 3582 1168 3586 1172
rect 70 1158 74 1162
rect 1774 1158 1778 1162
rect 1870 1158 1874 1162
rect 2142 1158 2146 1162
rect 2326 1158 2330 1162
rect 2350 1158 2354 1162
rect 2478 1158 2482 1162
rect 2502 1158 2506 1162
rect 2950 1158 2954 1162
rect 3030 1158 3034 1162
rect 3198 1158 3202 1162
rect 3478 1158 3482 1162
rect 6 1148 10 1152
rect 870 1148 874 1152
rect 934 1148 938 1152
rect 1006 1148 1010 1152
rect 1318 1148 1322 1152
rect 1558 1148 1562 1152
rect 1678 1148 1682 1152
rect 1686 1148 1690 1152
rect 1766 1148 1770 1152
rect 2150 1148 2154 1152
rect 2302 1148 2306 1152
rect 2374 1148 2378 1152
rect 2430 1148 2434 1152
rect 2438 1148 2442 1152
rect 2678 1148 2682 1152
rect 2878 1148 2882 1152
rect 2966 1148 2970 1152
rect 3206 1148 3210 1152
rect 3318 1148 3322 1152
rect 3534 1148 3538 1152
rect 710 1138 714 1142
rect 1022 1138 1026 1142
rect 1038 1138 1042 1142
rect 1046 1138 1050 1142
rect 1078 1138 1082 1142
rect 1166 1138 1170 1142
rect 1254 1138 1258 1142
rect 1814 1138 1818 1142
rect 1966 1138 1970 1142
rect 2030 1138 2034 1142
rect 2214 1138 2218 1142
rect 3070 1138 3074 1142
rect 3278 1138 3282 1142
rect 3334 1138 3338 1142
rect 534 1128 538 1132
rect 1246 1128 1250 1132
rect 1262 1128 1266 1132
rect 1406 1128 1410 1132
rect 1422 1128 1426 1132
rect 1430 1128 1434 1132
rect 1518 1128 1522 1132
rect 1534 1128 1538 1132
rect 1542 1128 1546 1132
rect 1590 1128 1594 1132
rect 478 1118 482 1122
rect 1950 1128 1954 1132
rect 2486 1128 2490 1132
rect 2558 1128 2562 1132
rect 2670 1128 2674 1132
rect 2726 1128 2730 1132
rect 2750 1128 2754 1132
rect 2998 1128 3002 1132
rect 3046 1128 3050 1132
rect 3126 1128 3130 1132
rect 3134 1128 3138 1132
rect 3190 1128 3194 1132
rect 3390 1128 3394 1132
rect 1102 1118 1106 1122
rect 1246 1118 1250 1122
rect 1382 1118 1386 1122
rect 1478 1118 1482 1122
rect 1598 1118 1602 1122
rect 1638 1118 1642 1122
rect 1854 1118 1858 1122
rect 2046 1118 2050 1122
rect 2118 1118 2122 1122
rect 2174 1118 2178 1122
rect 2470 1118 2474 1122
rect 2486 1118 2490 1122
rect 2598 1118 2602 1122
rect 2614 1118 2618 1122
rect 2662 1118 2666 1122
rect 2958 1118 2962 1122
rect 3198 1118 3202 1122
rect 3214 1118 3218 1122
rect 3422 1118 3426 1122
rect 3510 1118 3514 1122
rect 3630 1118 3634 1122
rect 830 1108 834 1112
rect 1270 1108 1274 1112
rect 1870 1108 1874 1112
rect 2166 1108 2170 1112
rect 2942 1108 2946 1112
rect 3110 1108 3114 1112
rect 3590 1108 3594 1112
rect 850 1103 854 1107
rect 858 1103 861 1107
rect 861 1103 862 1107
rect 1882 1103 1886 1107
rect 1890 1103 1893 1107
rect 1893 1103 1894 1107
rect 2906 1103 2910 1107
rect 2914 1103 2917 1107
rect 2917 1103 2918 1107
rect 366 1098 370 1102
rect 430 1098 434 1102
rect 966 1098 970 1102
rect 2934 1098 2938 1102
rect 3022 1098 3026 1102
rect 3462 1098 3466 1102
rect 3646 1098 3650 1102
rect 838 1088 842 1092
rect 1566 1088 1570 1092
rect 2126 1088 2130 1092
rect 158 1078 162 1082
rect 238 1078 242 1082
rect 1118 1078 1122 1082
rect 1158 1078 1162 1082
rect 1214 1078 1218 1082
rect 1238 1078 1242 1082
rect 1318 1078 1322 1082
rect 1662 1078 1666 1082
rect 1678 1078 1682 1082
rect 1766 1078 1770 1082
rect 1902 1078 1906 1082
rect 1958 1078 1962 1082
rect 2054 1078 2058 1082
rect 2670 1088 2674 1092
rect 2694 1088 2698 1092
rect 2750 1088 2754 1092
rect 3014 1088 3018 1092
rect 3094 1088 3098 1092
rect 3190 1088 3194 1092
rect 3246 1088 3250 1092
rect 3326 1088 3330 1092
rect 2086 1078 2090 1082
rect 2206 1078 2210 1082
rect 2326 1078 2330 1082
rect 2502 1078 2506 1082
rect 2518 1078 2522 1082
rect 2606 1078 2610 1082
rect 2646 1078 2650 1082
rect 3502 1078 3506 1082
rect 3526 1078 3530 1082
rect 3606 1078 3610 1082
rect 550 1068 554 1072
rect 902 1068 906 1072
rect 974 1068 978 1072
rect 1342 1068 1346 1072
rect 1558 1068 1562 1072
rect 1646 1068 1650 1072
rect 1934 1068 1938 1072
rect 2182 1068 2186 1072
rect 2430 1068 2434 1072
rect 2478 1068 2482 1072
rect 2670 1068 2674 1072
rect 2758 1068 2762 1072
rect 2814 1068 2818 1072
rect 2854 1068 2858 1072
rect 2862 1068 2866 1072
rect 3350 1068 3354 1072
rect 3422 1068 3426 1072
rect 3462 1068 3466 1072
rect 3486 1068 3490 1072
rect 3550 1068 3554 1072
rect 3710 1068 3714 1072
rect 22 1058 26 1062
rect 46 1058 50 1062
rect 334 1058 338 1062
rect 942 1058 946 1062
rect 998 1058 1002 1062
rect 1510 1058 1514 1062
rect 1526 1058 1530 1062
rect 2174 1058 2178 1062
rect 2190 1058 2194 1062
rect 2454 1058 2458 1062
rect 2486 1058 2490 1062
rect 2558 1058 2562 1062
rect 2574 1058 2578 1062
rect 2606 1058 2610 1062
rect 2638 1058 2642 1062
rect 2806 1058 2810 1062
rect 2886 1058 2890 1062
rect 3046 1058 3050 1062
rect 3070 1058 3074 1062
rect 3198 1058 3202 1062
rect 3286 1058 3290 1062
rect 3302 1058 3306 1062
rect 3526 1058 3530 1062
rect 3558 1058 3562 1062
rect 3614 1058 3618 1062
rect 678 1048 682 1052
rect 1358 1048 1362 1052
rect 1406 1048 1410 1052
rect 1422 1048 1426 1052
rect 1654 1048 1658 1052
rect 1662 1048 1666 1052
rect 1774 1048 1778 1052
rect 2102 1048 2106 1052
rect 2118 1048 2122 1052
rect 2438 1048 2442 1052
rect 2630 1048 2634 1052
rect 2710 1048 2714 1052
rect 2750 1048 2754 1052
rect 2830 1048 2834 1052
rect 3102 1048 3106 1052
rect 3454 1048 3458 1052
rect 3486 1048 3490 1052
rect 3510 1048 3514 1052
rect 486 1038 490 1042
rect 886 1038 890 1042
rect 1422 1038 1426 1042
rect 1494 1038 1498 1042
rect 1990 1038 1994 1042
rect 2558 1038 2562 1042
rect 2870 1038 2874 1042
rect 3478 1038 3482 1042
rect 1150 1028 1154 1032
rect 1350 1028 1354 1032
rect 1766 1028 1770 1032
rect 1838 1028 1842 1032
rect 2838 1028 2842 1032
rect 3166 1028 3170 1032
rect 3222 1028 3226 1032
rect 3510 1028 3514 1032
rect 3606 1028 3610 1032
rect 1102 1018 1106 1022
rect 1718 1018 1722 1022
rect 3030 1018 3034 1022
rect 3038 1018 3042 1022
rect 3046 1018 3050 1022
rect 3710 1018 3714 1022
rect 422 1008 426 1012
rect 1646 1008 1650 1012
rect 346 1003 350 1007
rect 354 1003 357 1007
rect 357 1003 358 1007
rect 1362 1003 1366 1007
rect 1370 1003 1373 1007
rect 1373 1003 1374 1007
rect 2386 1003 2390 1007
rect 2394 1003 2397 1007
rect 2397 1003 2398 1007
rect 3410 1003 3414 1007
rect 3418 1003 3421 1007
rect 3421 1003 3422 1007
rect 1254 998 1258 1002
rect 1582 998 1586 1002
rect 1670 998 1674 1002
rect 2182 998 2186 1002
rect 2566 998 2570 1002
rect 2934 998 2938 1002
rect 3070 998 3074 1002
rect 3166 998 3170 1002
rect 3638 998 3642 1002
rect 390 988 394 992
rect 3294 988 3298 992
rect 2118 978 2122 982
rect 2158 978 2162 982
rect 2574 978 2578 982
rect 2990 978 2994 982
rect 3030 978 3034 982
rect 3142 978 3146 982
rect 334 968 338 972
rect 958 968 962 972
rect 1854 968 1858 972
rect 1958 968 1962 972
rect 1966 968 1970 972
rect 2598 968 2602 972
rect 2926 968 2930 972
rect 2950 968 2954 972
rect 3086 968 3090 972
rect 3158 968 3162 972
rect 3230 968 3234 972
rect 3566 968 3570 972
rect 478 958 482 962
rect 646 958 650 962
rect 1606 958 1610 962
rect 1622 958 1626 962
rect 1718 958 1722 962
rect 1974 958 1978 962
rect 2390 958 2394 962
rect 2534 958 2538 962
rect 2558 958 2562 962
rect 2566 958 2570 962
rect 2686 958 2690 962
rect 2718 958 2722 962
rect 2830 958 2834 962
rect 2846 958 2850 962
rect 3150 958 3154 962
rect 3246 958 3250 962
rect 3366 958 3370 962
rect 3478 958 3482 962
rect 3486 958 3490 962
rect 310 948 314 952
rect 470 948 474 952
rect 1550 948 1554 952
rect 1726 948 1730 952
rect 1822 948 1826 952
rect 1910 948 1914 952
rect 1918 948 1922 952
rect 2166 948 2170 952
rect 2278 948 2282 952
rect 2286 948 2290 952
rect 2342 948 2346 952
rect 2366 948 2370 952
rect 2374 948 2378 952
rect 2414 948 2418 952
rect 2526 948 2530 952
rect 2582 948 2586 952
rect 2630 948 2634 952
rect 2662 948 2666 952
rect 2702 948 2706 952
rect 2742 948 2746 952
rect 2766 948 2770 952
rect 2806 948 2810 952
rect 2838 948 2842 952
rect 2870 948 2874 952
rect 2966 948 2970 952
rect 2974 948 2978 952
rect 2998 948 3002 952
rect 3062 948 3066 952
rect 3126 948 3130 952
rect 3254 948 3258 952
rect 3542 958 3546 962
rect 3630 958 3634 962
rect 3510 948 3514 952
rect 3526 948 3530 952
rect 286 938 290 942
rect 670 938 674 942
rect 790 938 794 942
rect 830 938 834 942
rect 1006 938 1010 942
rect 1542 938 1546 942
rect 1566 938 1570 942
rect 1590 938 1594 942
rect 1814 938 1818 942
rect 1846 938 1850 942
rect 2054 938 2058 942
rect 2534 938 2538 942
rect 2662 938 2666 942
rect 2678 938 2682 942
rect 2686 938 2690 942
rect 2742 938 2746 942
rect 3006 938 3010 942
rect 3062 938 3066 942
rect 3190 938 3194 942
rect 3270 938 3274 942
rect 3486 938 3490 942
rect 3566 938 3570 942
rect 334 928 338 932
rect 406 928 410 932
rect 598 928 602 932
rect 1046 928 1050 932
rect 1710 928 1714 932
rect 2198 928 2202 932
rect 2390 928 2394 932
rect 2622 928 2626 932
rect 2646 928 2650 932
rect 2862 928 2866 932
rect 2966 928 2970 932
rect 3182 928 3186 932
rect 3270 928 3274 932
rect 3510 928 3514 932
rect 422 918 426 922
rect 1726 918 1730 922
rect 2630 918 2634 922
rect 3358 918 3362 922
rect 3670 918 3674 922
rect 126 908 130 912
rect 822 908 826 912
rect 1798 908 1802 912
rect 2062 908 2066 912
rect 2078 908 2082 912
rect 2190 908 2194 912
rect 2414 908 2418 912
rect 2582 908 2586 912
rect 2710 908 2714 912
rect 2894 908 2898 912
rect 3662 908 3666 912
rect 850 903 854 907
rect 858 903 861 907
rect 861 903 862 907
rect 1882 903 1886 907
rect 1890 903 1893 907
rect 1893 903 1894 907
rect 2906 903 2910 907
rect 2914 903 2917 907
rect 2917 903 2918 907
rect 174 898 178 902
rect 1110 898 1114 902
rect 1590 898 1594 902
rect 1638 898 1642 902
rect 1846 898 1850 902
rect 2614 898 2618 902
rect 2766 898 2770 902
rect 2870 898 2874 902
rect 3030 898 3034 902
rect 3294 898 3298 902
rect 318 888 322 892
rect 406 888 410 892
rect 430 888 434 892
rect 462 888 466 892
rect 958 888 962 892
rect 1318 888 1322 892
rect 1894 888 1898 892
rect 1958 888 1962 892
rect 2254 888 2258 892
rect 3094 888 3098 892
rect 86 878 90 882
rect 206 878 210 882
rect 574 878 578 882
rect 686 878 690 882
rect 1006 878 1010 882
rect 1118 878 1122 882
rect 1286 878 1290 882
rect 1310 878 1314 882
rect 1454 878 1458 882
rect 1558 878 1562 882
rect 1766 878 1770 882
rect 1910 878 1914 882
rect 2374 878 2378 882
rect 2422 878 2426 882
rect 2502 878 2506 882
rect 2830 878 2834 882
rect 2854 878 2858 882
rect 2878 878 2882 882
rect 3070 878 3074 882
rect 3086 878 3090 882
rect 3294 878 3298 882
rect 3302 878 3306 882
rect 3326 878 3330 882
rect 3382 878 3386 882
rect 3406 878 3410 882
rect 3446 878 3450 882
rect 502 868 506 872
rect 646 868 650 872
rect 1022 868 1026 872
rect 1094 868 1098 872
rect 1142 868 1146 872
rect 1278 868 1282 872
rect 1486 868 1490 872
rect 1502 868 1506 872
rect 1774 868 1778 872
rect 1974 868 1978 872
rect 2054 868 2058 872
rect 2502 868 2506 872
rect 2518 868 2522 872
rect 2622 868 2626 872
rect 2678 868 2682 872
rect 2750 868 2754 872
rect 2814 868 2818 872
rect 2846 868 2850 872
rect 2854 868 2858 872
rect 2910 868 2914 872
rect 2918 868 2922 872
rect 2950 868 2954 872
rect 2974 868 2978 872
rect 3006 868 3010 872
rect 3158 868 3162 872
rect 3590 868 3594 872
rect 3622 868 3626 872
rect 374 858 378 862
rect 1126 858 1130 862
rect 1134 858 1138 862
rect 1350 858 1354 862
rect 1870 858 1874 862
rect 1966 858 1970 862
rect 2430 858 2434 862
rect 2694 858 2698 862
rect 2774 858 2778 862
rect 2790 858 2794 862
rect 3102 858 3106 862
rect 3206 858 3210 862
rect 3694 858 3698 862
rect 1414 848 1418 852
rect 1566 848 1570 852
rect 1814 848 1818 852
rect 1830 848 1834 852
rect 2030 848 2034 852
rect 2406 848 2410 852
rect 2654 848 2658 852
rect 2958 848 2962 852
rect 3478 848 3482 852
rect 3638 848 3642 852
rect 1150 838 1154 842
rect 1982 838 1986 842
rect 2902 838 2906 842
rect 2982 838 2986 842
rect 3006 838 3010 842
rect 3262 838 3266 842
rect 38 828 42 832
rect 1398 828 1402 832
rect 1934 828 1938 832
rect 1942 828 1946 832
rect 1950 828 1954 832
rect 2534 828 2538 832
rect 3070 828 3074 832
rect 3646 828 3650 832
rect 3686 828 3690 832
rect 166 818 170 822
rect 662 818 666 822
rect 734 818 738 822
rect 1294 818 1298 822
rect 1310 818 1314 822
rect 2118 818 2122 822
rect 2134 818 2138 822
rect 2798 818 2802 822
rect 3038 818 3042 822
rect 3142 818 3146 822
rect 3486 818 3490 822
rect 1630 808 1634 812
rect 2222 808 2226 812
rect 2454 808 2458 812
rect 2486 808 2490 812
rect 3182 808 3186 812
rect 3454 808 3458 812
rect 346 803 350 807
rect 354 803 357 807
rect 357 803 358 807
rect 1362 803 1366 807
rect 1370 803 1373 807
rect 1373 803 1374 807
rect 2386 803 2390 807
rect 2394 803 2397 807
rect 2397 803 2398 807
rect 3410 803 3414 807
rect 3418 803 3421 807
rect 3421 803 3422 807
rect 1854 798 1858 802
rect 1870 798 1874 802
rect 2150 798 2154 802
rect 2182 798 2186 802
rect 2494 798 2498 802
rect 3222 798 3226 802
rect 3606 798 3610 802
rect 2838 788 2842 792
rect 2982 788 2986 792
rect 3662 788 3666 792
rect 270 778 274 782
rect 806 778 810 782
rect 1166 778 1170 782
rect 2150 778 2154 782
rect 2182 778 2186 782
rect 2222 778 2226 782
rect 2286 778 2290 782
rect 2342 778 2346 782
rect 2462 778 2466 782
rect 2702 778 2706 782
rect 3014 778 3018 782
rect 3230 778 3234 782
rect 3366 778 3370 782
rect 3590 778 3594 782
rect 398 768 402 772
rect 886 768 890 772
rect 1510 768 1514 772
rect 2294 768 2298 772
rect 2302 768 2306 772
rect 2422 768 2426 772
rect 2766 768 2770 772
rect 2966 768 2970 772
rect 3014 768 3018 772
rect 3054 768 3058 772
rect 3590 768 3594 772
rect 310 758 314 762
rect 678 760 682 762
rect 678 758 682 760
rect 838 758 842 762
rect 1310 758 1314 762
rect 1542 758 1546 762
rect 1574 758 1578 762
rect 1766 758 1770 762
rect 1806 758 1810 762
rect 2582 758 2586 762
rect 2622 758 2626 762
rect 2830 758 2834 762
rect 2902 758 2906 762
rect 3254 758 3258 762
rect 3446 758 3450 762
rect 3542 758 3546 762
rect 3774 758 3778 762
rect 70 748 74 752
rect 238 748 242 752
rect 790 748 794 752
rect 1510 748 1514 752
rect 1566 748 1570 752
rect 1750 748 1754 752
rect 2262 748 2266 752
rect 2430 748 2434 752
rect 2494 748 2498 752
rect 2518 748 2522 752
rect 2686 748 2690 752
rect 2702 748 2706 752
rect 1814 738 1818 742
rect 1950 738 1954 742
rect 2854 748 2858 752
rect 2926 748 2930 752
rect 2990 748 2994 752
rect 3054 748 3058 752
rect 3598 748 3602 752
rect 2486 738 2490 742
rect 2982 738 2986 742
rect 3206 738 3210 742
rect 3246 738 3250 742
rect 3302 738 3306 742
rect 3574 738 3578 742
rect 622 728 626 732
rect 654 728 658 732
rect 1006 728 1010 732
rect 1150 728 1154 732
rect 1710 728 1714 732
rect 1998 728 2002 732
rect 2382 728 2386 732
rect 2478 728 2482 732
rect 2630 728 2634 732
rect 2678 728 2682 732
rect 2686 728 2690 732
rect 2894 728 2898 732
rect 2950 728 2954 732
rect 3046 728 3050 732
rect 3062 728 3066 732
rect 3110 728 3114 732
rect 3294 728 3298 732
rect 102 718 106 722
rect 750 718 754 722
rect 3454 728 3458 732
rect 3462 728 3466 732
rect 3622 728 3626 732
rect 3710 728 3714 732
rect 1510 718 1514 722
rect 3078 718 3082 722
rect 3182 718 3186 722
rect 3318 718 3322 722
rect 3334 718 3338 722
rect 3374 718 3378 722
rect 3614 718 3618 722
rect 3670 718 3674 722
rect 590 708 594 712
rect 1118 708 1122 712
rect 1918 708 1922 712
rect 2406 708 2410 712
rect 2862 708 2866 712
rect 2926 708 2930 712
rect 3318 708 3322 712
rect 3598 708 3602 712
rect 3678 708 3682 712
rect 850 703 854 707
rect 858 703 861 707
rect 861 703 862 707
rect 1882 703 1886 707
rect 1890 703 1893 707
rect 1893 703 1894 707
rect 2906 703 2910 707
rect 2914 703 2917 707
rect 2917 703 2918 707
rect 166 698 170 702
rect 662 698 666 702
rect 2174 698 2178 702
rect 2822 698 2826 702
rect 2854 698 2858 702
rect 3294 698 3298 702
rect 3558 698 3562 702
rect 3622 698 3626 702
rect 3758 698 3762 702
rect 1046 688 1050 692
rect 1598 688 1602 692
rect 2254 688 2258 692
rect 2294 688 2298 692
rect 2470 688 2474 692
rect 2478 688 2482 692
rect 2774 688 2778 692
rect 2806 688 2810 692
rect 2998 688 3002 692
rect 3294 688 3298 692
rect 3622 688 3626 692
rect 86 678 90 682
rect 414 678 418 682
rect 494 678 498 682
rect 1150 678 1154 682
rect 1462 678 1466 682
rect 1494 678 1498 682
rect 1742 678 1746 682
rect 1966 678 1970 682
rect 2262 678 2266 682
rect 2446 678 2450 682
rect 2502 678 2506 682
rect 2870 678 2874 682
rect 3006 678 3010 682
rect 3366 678 3370 682
rect 3398 678 3402 682
rect 3502 678 3506 682
rect 374 668 378 672
rect 422 668 426 672
rect 526 668 530 672
rect 582 668 586 672
rect 638 668 642 672
rect 1422 668 1426 672
rect 1598 668 1602 672
rect 1950 668 1954 672
rect 1958 668 1962 672
rect 2278 668 2282 672
rect 2470 668 2474 672
rect 2782 668 2786 672
rect 3094 668 3098 672
rect 3278 668 3282 672
rect 214 658 218 662
rect 398 658 402 662
rect 1246 658 1250 662
rect 1654 658 1658 662
rect 1926 658 1930 662
rect 2038 658 2042 662
rect 2102 658 2106 662
rect 2174 658 2178 662
rect 2342 658 2346 662
rect 2662 658 2666 662
rect 2998 658 3002 662
rect 3038 658 3042 662
rect 3118 658 3122 662
rect 3166 658 3170 662
rect 3206 658 3210 662
rect 3590 658 3594 662
rect 3670 658 3674 662
rect 1454 648 1458 652
rect 1726 648 1730 652
rect 1998 648 2002 652
rect 2006 648 2010 652
rect 2366 648 2370 652
rect 2494 648 2498 652
rect 2582 648 2586 652
rect 3174 648 3178 652
rect 3558 648 3562 652
rect 3758 648 3762 652
rect 2246 638 2250 642
rect 2318 638 2322 642
rect 2774 638 2778 642
rect 2790 638 2794 642
rect 2798 638 2802 642
rect 2878 638 2882 642
rect 2902 638 2906 642
rect 3254 638 3258 642
rect 3678 638 3682 642
rect 1278 628 1282 632
rect 1710 628 1714 632
rect 1942 628 1946 632
rect 2254 628 2258 632
rect 3102 628 3106 632
rect 3382 628 3386 632
rect 1838 618 1842 622
rect 2366 618 2370 622
rect 2374 618 2378 622
rect 3510 618 3514 622
rect 870 608 874 612
rect 2014 608 2018 612
rect 2022 608 2026 612
rect 2206 608 2210 612
rect 2766 608 2770 612
rect 2774 608 2778 612
rect 3310 608 3314 612
rect 3430 608 3434 612
rect 346 603 350 607
rect 354 603 357 607
rect 357 603 358 607
rect 1362 603 1366 607
rect 1370 603 1373 607
rect 1373 603 1374 607
rect 2386 603 2390 607
rect 2394 603 2397 607
rect 2397 603 2398 607
rect 3410 603 3414 607
rect 3418 603 3421 607
rect 3421 603 3422 607
rect 1454 598 1458 602
rect 2086 598 2090 602
rect 2094 598 2098 602
rect 2142 598 2146 602
rect 2486 598 2490 602
rect 2534 598 2538 602
rect 2718 598 2722 602
rect 3118 598 3122 602
rect 3670 598 3674 602
rect 1390 588 1394 592
rect 1598 588 1602 592
rect 2070 588 2074 592
rect 2366 588 2370 592
rect 2374 588 2378 592
rect 2526 588 2530 592
rect 2726 588 2730 592
rect 3454 588 3458 592
rect 230 578 234 582
rect 974 578 978 582
rect 1534 578 1538 582
rect 1718 578 1722 582
rect 3118 578 3122 582
rect 3670 578 3674 582
rect 782 568 786 572
rect 1142 568 1146 572
rect 1246 568 1250 572
rect 1406 568 1410 572
rect 2822 568 2826 572
rect 2926 568 2930 572
rect 2934 568 2938 572
rect 2998 568 3002 572
rect 238 558 242 562
rect 366 558 370 562
rect 1646 558 1650 562
rect 2158 558 2162 562
rect 2230 558 2234 562
rect 2302 558 2306 562
rect 2334 558 2338 562
rect 2694 558 2698 562
rect 2846 558 2850 562
rect 2854 558 2858 562
rect 2958 558 2962 562
rect 3158 558 3162 562
rect 3190 558 3194 562
rect 3214 558 3218 562
rect 3598 558 3602 562
rect 1318 548 1322 552
rect 1390 548 1394 552
rect 1438 548 1442 552
rect 1614 548 1618 552
rect 2590 548 2594 552
rect 2710 548 2714 552
rect 2934 548 2938 552
rect 3174 548 3178 552
rect 3206 548 3210 552
rect 3430 548 3434 552
rect 3502 548 3506 552
rect 3550 548 3554 552
rect 270 538 274 542
rect 902 538 906 542
rect 1030 538 1034 542
rect 1110 538 1114 542
rect 1366 538 1370 542
rect 1446 538 1450 542
rect 1950 538 1954 542
rect 2518 538 2522 542
rect 2622 538 2626 542
rect 2742 538 2746 542
rect 2806 538 2810 542
rect 3078 538 3082 542
rect 3462 538 3466 542
rect 3510 538 3514 542
rect 3558 538 3562 542
rect 382 528 386 532
rect 1246 528 1250 532
rect 1550 528 1554 532
rect 1614 528 1618 532
rect 1790 528 1794 532
rect 2350 528 2354 532
rect 2454 528 2458 532
rect 2926 528 2930 532
rect 3278 528 3282 532
rect 3414 528 3418 532
rect 3486 528 3490 532
rect 3710 528 3714 532
rect 62 518 66 522
rect 1574 518 1578 522
rect 1590 518 1594 522
rect 2134 518 2138 522
rect 2774 518 2778 522
rect 2806 518 2810 522
rect 142 508 146 512
rect 1278 508 1282 512
rect 1438 508 1442 512
rect 1558 508 1562 512
rect 2894 508 2898 512
rect 3286 508 3290 512
rect 3510 508 3514 512
rect 850 503 854 507
rect 858 503 861 507
rect 861 503 862 507
rect 1882 503 1886 507
rect 1890 503 1893 507
rect 1893 503 1894 507
rect 2906 503 2910 507
rect 2914 503 2917 507
rect 2917 503 2918 507
rect 70 498 74 502
rect 1382 498 1386 502
rect 1438 498 1442 502
rect 1446 498 1450 502
rect 1718 498 1722 502
rect 1726 498 1730 502
rect 2054 498 2058 502
rect 2446 498 2450 502
rect 2862 498 2866 502
rect 2926 498 2930 502
rect 3270 498 3274 502
rect 3654 498 3658 502
rect 3718 498 3722 502
rect 798 488 802 492
rect 1014 488 1018 492
rect 1590 488 1594 492
rect 1854 488 1858 492
rect 2094 488 2098 492
rect 2790 488 2794 492
rect 2814 488 2818 492
rect 2862 488 2866 492
rect 3102 488 3106 492
rect 3342 488 3346 492
rect 3542 488 3546 492
rect 86 478 90 482
rect 806 478 810 482
rect 1534 478 1538 482
rect 1606 478 1610 482
rect 1798 478 1802 482
rect 1846 478 1850 482
rect 2214 478 2218 482
rect 2382 478 2386 482
rect 2446 478 2450 482
rect 2470 478 2474 482
rect 2494 478 2498 482
rect 2590 478 2594 482
rect 2838 478 2842 482
rect 3222 478 3226 482
rect 3454 478 3458 482
rect 3558 478 3562 482
rect 3654 478 3658 482
rect 870 468 874 472
rect 1390 468 1394 472
rect 1750 468 1754 472
rect 1814 468 1818 472
rect 1822 468 1826 472
rect 1934 468 1938 472
rect 1950 468 1954 472
rect 2110 468 2114 472
rect 2182 468 2186 472
rect 2558 468 2562 472
rect 2654 468 2658 472
rect 2854 468 2858 472
rect 222 458 226 462
rect 1246 458 1250 462
rect 1286 458 1290 462
rect 1382 458 1386 462
rect 1430 458 1434 462
rect 1446 458 1450 462
rect 1558 458 1562 462
rect 2246 458 2250 462
rect 2318 458 2322 462
rect 2382 458 2386 462
rect 2486 458 2490 462
rect 2718 458 2722 462
rect 2742 458 2746 462
rect 2870 458 2874 462
rect 2934 458 2938 462
rect 2958 458 2962 462
rect 2982 458 2986 462
rect 3430 458 3434 462
rect 3574 458 3578 462
rect 3702 458 3706 462
rect 838 448 842 452
rect 926 448 930 452
rect 1518 448 1522 452
rect 1598 448 1602 452
rect 1974 448 1978 452
rect 2550 448 2554 452
rect 2854 448 2858 452
rect 3038 448 3042 452
rect 3214 448 3218 452
rect 3302 448 3306 452
rect 3574 448 3578 452
rect 3670 448 3674 452
rect 1158 438 1162 442
rect 1230 438 1234 442
rect 1486 438 1490 442
rect 1542 438 1546 442
rect 2086 438 2090 442
rect 2366 438 2370 442
rect 2374 438 2378 442
rect 2486 438 2490 442
rect 2622 438 2626 442
rect 2694 438 2698 442
rect 3518 438 3522 442
rect 558 428 562 432
rect 2030 428 2034 432
rect 2574 428 2578 432
rect 2646 428 2650 432
rect 2790 428 2794 432
rect 3022 428 3026 432
rect 3134 428 3138 432
rect 902 418 906 422
rect 1262 418 1266 422
rect 2238 418 2242 422
rect 2342 418 2346 422
rect 3174 418 3178 422
rect 622 408 626 412
rect 1406 408 1410 412
rect 1814 408 1818 412
rect 2854 408 2858 412
rect 2878 408 2882 412
rect 3534 408 3538 412
rect 346 403 350 407
rect 354 403 357 407
rect 357 403 358 407
rect 1362 403 1366 407
rect 1370 403 1373 407
rect 1373 403 1374 407
rect 2386 403 2390 407
rect 2394 403 2397 407
rect 2397 403 2398 407
rect 3410 403 3414 407
rect 3418 403 3421 407
rect 3421 403 3422 407
rect 1350 398 1354 402
rect 1582 398 1586 402
rect 2542 398 2546 402
rect 2790 398 2794 402
rect 2966 398 2970 402
rect 3022 398 3026 402
rect 582 388 586 392
rect 1078 388 1082 392
rect 2134 388 2138 392
rect 2190 388 2194 392
rect 2398 388 2402 392
rect 2430 388 2434 392
rect 2630 388 2634 392
rect 3014 388 3018 392
rect 974 378 978 382
rect 1350 378 1354 382
rect 2038 378 2042 382
rect 2046 378 2050 382
rect 2094 378 2098 382
rect 2142 378 2146 382
rect 2246 378 2250 382
rect 2526 378 2530 382
rect 2742 378 2746 382
rect 2990 378 2994 382
rect 1110 368 1114 372
rect 1942 368 1946 372
rect 2510 368 2514 372
rect 3150 368 3154 372
rect 3638 368 3642 372
rect 310 358 314 362
rect 1686 358 1690 362
rect 1838 358 1842 362
rect 2014 358 2018 362
rect 2246 358 2250 362
rect 2310 358 2314 362
rect 2374 358 2378 362
rect 2750 358 2754 362
rect 3158 358 3162 362
rect 3214 358 3218 362
rect 3454 358 3458 362
rect 3638 358 3642 362
rect 3670 358 3674 362
rect 590 348 594 352
rect 974 348 978 352
rect 1110 348 1114 352
rect 1142 348 1146 352
rect 1862 348 1866 352
rect 1950 348 1954 352
rect 2326 348 2330 352
rect 2350 348 2354 352
rect 2494 348 2498 352
rect 2566 348 2570 352
rect 2702 348 2706 352
rect 2726 348 2730 352
rect 2734 348 2738 352
rect 2846 348 2850 352
rect 2870 348 2874 352
rect 2926 348 2930 352
rect 3014 348 3018 352
rect 3558 348 3562 352
rect 3662 348 3666 352
rect 142 338 146 342
rect 534 338 538 342
rect 942 338 946 342
rect 1014 338 1018 342
rect 1390 338 1394 342
rect 1542 338 1546 342
rect 1838 338 1842 342
rect 1974 338 1978 342
rect 2046 338 2050 342
rect 2086 338 2090 342
rect 2270 338 2274 342
rect 2286 338 2290 342
rect 2334 338 2338 342
rect 2414 338 2418 342
rect 2462 338 2466 342
rect 2598 338 2602 342
rect 2750 338 2754 342
rect 2790 338 2794 342
rect 2854 338 2858 342
rect 3062 338 3066 342
rect 3222 338 3226 342
rect 3710 338 3714 342
rect 3758 338 3762 342
rect 734 328 738 332
rect 1094 328 1098 332
rect 1110 328 1114 332
rect 1742 328 1746 332
rect 2022 328 2026 332
rect 2230 328 2234 332
rect 2534 328 2538 332
rect 2654 328 2658 332
rect 2830 328 2834 332
rect 2894 328 2898 332
rect 3278 328 3282 332
rect 3518 328 3522 332
rect 3598 328 3602 332
rect 3622 328 3626 332
rect 3822 328 3826 332
rect 2710 318 2714 322
rect 2838 318 2842 322
rect 3174 318 3178 322
rect 3270 318 3274 322
rect 1870 308 1874 312
rect 2574 308 2578 312
rect 3030 308 3034 312
rect 850 303 854 307
rect 858 303 861 307
rect 861 303 862 307
rect 1882 303 1886 307
rect 1890 303 1893 307
rect 1893 303 1894 307
rect 2906 303 2910 307
rect 2914 303 2917 307
rect 2917 303 2918 307
rect 2470 298 2474 302
rect 2478 298 2482 302
rect 2590 298 2594 302
rect 2806 298 2810 302
rect 2894 298 2898 302
rect 2982 298 2986 302
rect 3470 298 3474 302
rect 494 288 498 292
rect 1094 288 1098 292
rect 1502 288 1506 292
rect 1622 288 1626 292
rect 1934 288 1938 292
rect 2030 288 2034 292
rect 2062 288 2066 292
rect 2150 288 2154 292
rect 2206 288 2210 292
rect 2222 288 2226 292
rect 2446 288 2450 292
rect 814 278 818 282
rect 1022 278 1026 282
rect 1294 278 1298 282
rect 1510 278 1514 282
rect 2054 278 2058 282
rect 2118 278 2122 282
rect 2134 278 2138 282
rect 2198 278 2202 282
rect 2214 278 2218 282
rect 2230 278 2234 282
rect 2310 278 2314 282
rect 2870 278 2874 282
rect 3126 278 3130 282
rect 3190 278 3194 282
rect 3342 278 3346 282
rect 70 268 74 272
rect 286 268 290 272
rect 478 268 482 272
rect 550 268 554 272
rect 1102 268 1106 272
rect 1382 268 1386 272
rect 1518 268 1522 272
rect 1534 268 1538 272
rect 1574 268 1578 272
rect 1590 268 1594 272
rect 1614 268 1618 272
rect 1750 268 1754 272
rect 2598 268 2602 272
rect 2606 268 2610 272
rect 2862 268 2866 272
rect 3350 268 3354 272
rect 3574 268 3578 272
rect 3614 268 3618 272
rect 558 258 562 262
rect 662 258 666 262
rect 1958 258 1962 262
rect 2870 258 2874 262
rect 3006 258 3010 262
rect 3150 258 3154 262
rect 3286 258 3290 262
rect 1102 248 1106 252
rect 1526 248 1530 252
rect 1614 248 1618 252
rect 1622 248 1626 252
rect 1710 248 1714 252
rect 1766 248 1770 252
rect 1782 248 1786 252
rect 1926 248 1930 252
rect 1974 248 1978 252
rect 2238 248 2242 252
rect 2510 248 2514 252
rect 2518 248 2522 252
rect 3022 248 3026 252
rect 1182 238 1186 242
rect 1438 238 1442 242
rect 1558 238 1562 242
rect 1846 238 1850 242
rect 1950 238 1954 242
rect 2190 238 2194 242
rect 2206 228 2210 232
rect 1646 218 1650 222
rect 2470 218 2474 222
rect 2478 218 2482 222
rect 2838 218 2842 222
rect 3294 218 3298 222
rect 3734 218 3738 222
rect 86 208 90 212
rect 1342 208 1346 212
rect 3446 208 3450 212
rect 346 203 350 207
rect 354 203 357 207
rect 357 203 358 207
rect 1362 203 1366 207
rect 1370 203 1373 207
rect 1373 203 1374 207
rect 2386 203 2390 207
rect 2394 203 2397 207
rect 2397 203 2398 207
rect 3410 203 3414 207
rect 3418 203 3421 207
rect 3421 203 3422 207
rect 1350 198 1354 202
rect 1622 198 1626 202
rect 2014 198 2018 202
rect 2214 198 2218 202
rect 2286 198 2290 202
rect 3566 198 3570 202
rect 2046 188 2050 192
rect 2422 188 2426 192
rect 2478 188 2482 192
rect 2814 188 2818 192
rect 2974 188 2978 192
rect 3078 188 3082 192
rect 1030 178 1034 182
rect 1614 178 1618 182
rect 1654 178 1658 182
rect 1662 178 1666 182
rect 1990 178 1994 182
rect 2926 178 2930 182
rect 3582 178 3586 182
rect 1286 168 1290 172
rect 1958 168 1962 172
rect 2174 168 2178 172
rect 2430 168 2434 172
rect 2710 168 2714 172
rect 3158 168 3162 172
rect 3550 168 3554 172
rect 3710 168 3714 172
rect 766 158 770 162
rect 1190 158 1194 162
rect 2230 158 2234 162
rect 2254 158 2258 162
rect 2686 158 2690 162
rect 2998 158 3002 162
rect 3574 158 3578 162
rect 38 148 42 152
rect 1214 148 1218 152
rect 1686 148 1690 152
rect 2142 148 2146 152
rect 2718 148 2722 152
rect 2894 148 2898 152
rect 3166 148 3170 152
rect 3558 148 3562 152
rect 3606 148 3610 152
rect 3686 148 3690 152
rect 3718 148 3722 152
rect 598 138 602 142
rect 1238 138 1242 142
rect 1742 138 1746 142
rect 2150 138 2154 142
rect 2222 138 2226 142
rect 2238 138 2242 142
rect 2686 138 2690 142
rect 3014 138 3018 142
rect 3030 138 3034 142
rect 3294 138 3298 142
rect 3422 138 3426 142
rect 3678 138 3682 142
rect 1070 128 1074 132
rect 1462 128 1466 132
rect 2558 128 2562 132
rect 3494 128 3498 132
rect 3710 128 3714 132
rect 774 118 778 122
rect 3318 118 3322 122
rect 2486 108 2490 112
rect 3238 108 3242 112
rect 3358 108 3362 112
rect 3742 108 3746 112
rect 850 103 854 107
rect 858 103 861 107
rect 861 103 862 107
rect 1882 103 1886 107
rect 1890 103 1893 107
rect 1893 103 1894 107
rect 2906 103 2910 107
rect 2914 103 2917 107
rect 2917 103 2918 107
rect 726 98 730 102
rect 1790 98 1794 102
rect 3134 98 3138 102
rect 3142 98 3146 102
rect 766 88 770 92
rect 1310 88 1314 92
rect 1646 88 1650 92
rect 2102 88 2106 92
rect 2502 88 2506 92
rect 3430 88 3434 92
rect 3638 88 3642 92
rect 910 78 914 82
rect 1806 78 1810 82
rect 2254 78 2258 82
rect 3134 78 3138 82
rect 3334 78 3338 82
rect 3710 78 3714 82
rect 502 68 506 72
rect 750 68 754 72
rect 1118 68 1122 72
rect 2102 68 2106 72
rect 2206 68 2210 72
rect 2606 68 2610 72
rect 2742 68 2746 72
rect 3230 68 3234 72
rect 3350 68 3354 72
rect 3582 68 3586 72
rect 3694 68 3698 72
rect 3758 68 3762 72
rect 574 58 578 62
rect 2038 58 2042 62
rect 3318 58 3322 62
rect 3374 58 3378 62
rect 3390 58 3394 62
rect 3486 58 3490 62
rect 3526 58 3530 62
rect 3766 58 3770 62
rect 2854 48 2858 52
rect 3726 48 3730 52
rect 3326 38 3330 42
rect 3382 38 3386 42
rect 1342 28 1346 32
rect 2014 28 2018 32
rect 3646 28 3650 32
rect 1214 18 1218 22
rect 1278 18 1282 22
rect 1926 18 1930 22
rect 2094 18 2098 22
rect 734 8 738 12
rect 1086 8 1090 12
rect 2510 8 2514 12
rect 346 3 350 7
rect 354 3 357 7
rect 357 3 358 7
rect 1362 3 1366 7
rect 1370 3 1373 7
rect 1373 3 1374 7
rect 2386 3 2390 7
rect 2394 3 2397 7
rect 2397 3 2398 7
rect 3410 3 3414 7
rect 3418 3 3421 7
rect 3421 3 3422 7
<< metal4 >>
rect 344 3603 346 3607
rect 350 3603 353 3607
rect 358 3603 360 3607
rect 1360 3603 1362 3607
rect 1366 3603 1369 3607
rect 1374 3603 1376 3607
rect 2384 3603 2386 3607
rect 2390 3603 2393 3607
rect 2398 3603 2400 3607
rect 3408 3603 3410 3607
rect 3414 3603 3417 3607
rect 3422 3603 3424 3607
rect 426 3598 433 3601
rect 286 3518 294 3521
rect 6 3142 9 3458
rect 138 3268 142 3271
rect 38 2852 41 2858
rect 62 2462 65 2858
rect 110 2842 113 3238
rect 122 2848 126 2851
rect 30 2192 33 2278
rect 6 1952 9 1958
rect 10 1848 14 1851
rect 6 1662 9 1668
rect 6 1522 9 1548
rect 10 1338 14 1341
rect 38 1272 41 2268
rect 46 1942 49 1948
rect 54 1942 57 2068
rect 62 1952 65 2058
rect 110 1912 113 2838
rect 134 2742 137 2748
rect 130 2508 137 2511
rect 134 2492 137 2508
rect 142 2261 145 2578
rect 142 2258 150 2261
rect 134 2132 137 2138
rect 142 1922 145 2258
rect 158 2002 161 2548
rect 190 2442 193 2468
rect 198 2262 201 3458
rect 230 3072 233 3298
rect 214 2522 217 2798
rect 214 2442 217 2518
rect 206 2402 209 2418
rect 126 1732 129 1878
rect 134 1732 137 1738
rect 94 1632 97 1678
rect 114 1668 118 1671
rect 10 1168 14 1171
rect 10 1148 14 1151
rect 22 1062 25 1068
rect 38 832 41 1268
rect 50 1058 54 1061
rect 38 152 41 828
rect 70 752 73 1158
rect 86 882 89 888
rect 62 522 65 728
rect 86 682 89 688
rect 70 272 73 498
rect 94 481 97 1628
rect 126 912 129 1728
rect 158 1082 161 1998
rect 194 1938 198 1941
rect 166 1242 169 1418
rect 182 1362 185 1418
rect 174 1322 177 1338
rect 102 722 105 728
rect 166 702 169 818
rect 174 692 177 898
rect 210 878 217 881
rect 214 662 217 878
rect 90 478 97 481
rect 86 212 89 478
rect 142 342 145 508
rect 222 462 225 3058
rect 230 2882 233 3068
rect 238 3062 241 3388
rect 286 3272 289 3518
rect 430 3512 433 3598
rect 1506 3598 1513 3601
rect 344 3403 346 3407
rect 350 3403 353 3407
rect 358 3403 360 3407
rect 558 3402 561 3438
rect 446 3258 454 3261
rect 318 3192 321 3248
rect 344 3203 346 3207
rect 350 3203 353 3207
rect 358 3203 360 3207
rect 318 2942 321 3188
rect 344 3003 346 3007
rect 350 3003 353 3007
rect 358 3003 360 3007
rect 250 2848 254 2851
rect 334 2752 337 2898
rect 344 2803 346 2807
rect 350 2803 353 2807
rect 358 2803 360 2807
rect 230 2032 233 2068
rect 238 1672 241 2478
rect 238 1482 241 1668
rect 230 582 233 1168
rect 238 1082 241 1478
rect 262 1242 265 2098
rect 270 1872 273 1948
rect 286 1731 289 2218
rect 294 1752 297 2258
rect 286 1728 294 1731
rect 286 942 289 1728
rect 302 1352 305 1558
rect 310 952 313 1748
rect 334 1672 337 2658
rect 344 2603 346 2607
rect 350 2603 353 2607
rect 358 2603 360 2607
rect 366 2482 369 3028
rect 374 2642 377 2648
rect 344 2403 346 2407
rect 350 2403 353 2407
rect 358 2403 360 2407
rect 344 2203 346 2207
rect 350 2203 353 2207
rect 358 2203 360 2207
rect 344 2003 346 2007
rect 350 2003 353 2007
rect 358 2003 360 2007
rect 344 1803 346 1807
rect 350 1803 353 1807
rect 358 1803 360 1807
rect 366 1712 369 2128
rect 374 1732 377 2468
rect 382 1752 385 2528
rect 344 1603 346 1607
rect 350 1603 353 1607
rect 358 1603 360 1607
rect 344 1403 346 1407
rect 350 1403 353 1407
rect 358 1403 360 1407
rect 382 1372 385 1748
rect 422 1732 425 2188
rect 446 2142 449 3258
rect 502 3132 505 3318
rect 558 3252 561 3398
rect 510 3242 513 3248
rect 454 2352 457 2868
rect 502 2662 505 2668
rect 462 2512 465 2658
rect 474 2638 481 2641
rect 478 2632 481 2638
rect 454 1862 457 2038
rect 462 1742 465 2298
rect 390 1482 393 1688
rect 344 1203 346 1207
rect 350 1203 353 1207
rect 358 1203 360 1207
rect 330 1058 334 1061
rect 344 1003 346 1007
rect 350 1003 353 1007
rect 358 1003 360 1007
rect 334 932 337 968
rect 318 892 321 898
rect 344 803 346 807
rect 350 803 353 807
rect 358 803 360 807
rect 238 562 241 748
rect 270 542 273 778
rect 310 362 313 758
rect 344 603 346 607
rect 350 603 353 607
rect 358 603 360 607
rect 366 562 369 1098
rect 374 672 377 858
rect 382 532 385 1278
rect 390 661 393 988
rect 406 892 409 928
rect 398 888 406 891
rect 398 772 401 888
rect 414 682 417 1728
rect 422 1012 425 1468
rect 430 1182 433 1508
rect 438 1292 441 1728
rect 462 1542 465 1698
rect 470 1562 473 2048
rect 478 1932 481 1938
rect 494 1922 497 2378
rect 478 1742 481 1748
rect 502 1702 505 2338
rect 510 1872 513 3238
rect 550 2772 553 2938
rect 518 2151 521 2708
rect 538 2468 542 2471
rect 550 2182 553 2768
rect 518 2148 526 2151
rect 526 2142 529 2148
rect 526 1982 529 2138
rect 558 2052 561 3248
rect 574 3112 577 3178
rect 566 2842 569 3068
rect 574 2932 577 3108
rect 582 3082 585 3428
rect 566 1972 569 2738
rect 582 2652 585 3008
rect 590 2992 593 3248
rect 598 3042 601 3128
rect 598 3032 601 3038
rect 606 2951 609 3258
rect 606 2948 614 2951
rect 606 2692 609 2948
rect 598 2602 601 2688
rect 614 2242 617 2758
rect 638 2671 641 2738
rect 634 2668 641 2671
rect 646 2672 649 3068
rect 638 2482 641 2668
rect 646 2562 649 2568
rect 654 2562 657 2798
rect 662 2731 665 3038
rect 670 2992 673 3538
rect 678 3332 681 3478
rect 686 2928 694 2931
rect 686 2812 689 2928
rect 662 2728 670 2731
rect 670 2652 673 2728
rect 666 2558 670 2561
rect 682 2368 686 2371
rect 646 2352 649 2368
rect 462 1292 465 1528
rect 486 1448 494 1451
rect 422 672 425 918
rect 430 892 433 1098
rect 454 891 457 1168
rect 470 952 473 1348
rect 478 1322 481 1328
rect 486 1322 489 1448
rect 478 962 481 1118
rect 486 1042 489 1268
rect 454 888 462 891
rect 502 872 505 1678
rect 526 1642 529 1658
rect 518 1482 521 1628
rect 534 1622 537 1748
rect 510 1172 513 1388
rect 534 1362 537 1618
rect 542 1332 545 1718
rect 494 682 497 688
rect 390 658 398 661
rect 382 492 385 528
rect 344 403 346 407
rect 350 403 353 407
rect 358 403 360 407
rect 494 292 497 678
rect 526 672 529 1308
rect 534 1132 537 1138
rect 542 902 545 1328
rect 550 1072 553 1878
rect 566 1402 569 1838
rect 562 1338 566 1341
rect 574 1332 577 2178
rect 590 1452 593 1858
rect 610 1848 614 1851
rect 562 1168 566 1171
rect 538 338 542 341
rect 478 272 481 278
rect 550 272 553 1068
rect 570 878 574 881
rect 582 672 585 1398
rect 622 1232 625 1918
rect 630 1862 633 2048
rect 638 1952 641 2148
rect 646 1828 654 1831
rect 646 1502 649 1828
rect 658 1738 662 1741
rect 290 268 294 271
rect 558 262 561 428
rect 344 203 346 207
rect 350 203 353 207
rect 358 203 360 207
rect 506 68 510 71
rect 582 61 585 388
rect 590 352 593 708
rect 598 142 601 928
rect 622 412 625 728
rect 638 672 641 1198
rect 646 872 649 958
rect 654 732 657 1478
rect 662 1472 665 1678
rect 670 1542 673 1748
rect 678 1652 681 2348
rect 694 2332 697 2548
rect 686 1732 689 1948
rect 702 1882 705 3468
rect 734 3412 737 3548
rect 848 3503 850 3507
rect 854 3503 857 3507
rect 862 3503 864 3507
rect 870 3432 873 3508
rect 894 3472 897 3598
rect 906 3538 910 3541
rect 774 3342 777 3418
rect 758 3248 766 3251
rect 726 3142 729 3158
rect 742 3072 745 3238
rect 758 3132 761 3248
rect 710 2842 713 2968
rect 750 2932 753 2938
rect 758 2932 761 3118
rect 710 2152 713 2778
rect 726 2668 734 2671
rect 726 2662 729 2668
rect 730 2638 734 2641
rect 718 2562 721 2638
rect 718 2452 721 2558
rect 734 2462 737 2468
rect 750 2432 753 2928
rect 766 2872 769 2998
rect 762 2858 766 2861
rect 762 2768 766 2771
rect 762 2678 766 2681
rect 774 2642 777 3338
rect 848 3303 850 3307
rect 854 3303 857 3307
rect 862 3303 864 3307
rect 942 3282 945 3418
rect 950 3282 953 3328
rect 782 3082 785 3268
rect 782 2902 785 3078
rect 814 2872 817 3148
rect 848 3103 850 3107
rect 854 3103 857 3107
rect 862 3103 864 3107
rect 710 1942 713 2148
rect 666 1388 670 1391
rect 694 1322 697 1878
rect 718 1782 721 2098
rect 734 2022 737 2158
rect 742 2152 745 2358
rect 758 2252 761 2538
rect 766 2182 769 2568
rect 754 2158 761 2161
rect 730 1948 734 1951
rect 718 1512 721 1668
rect 726 1592 729 1858
rect 742 1572 745 1938
rect 750 1932 753 2138
rect 758 2012 761 2158
rect 750 1662 753 1788
rect 670 942 673 1298
rect 734 1292 737 1488
rect 750 1422 753 1608
rect 758 1392 761 1938
rect 774 1922 777 2638
rect 782 2522 785 2768
rect 790 2392 793 2868
rect 814 2792 817 2868
rect 806 2772 809 2778
rect 822 2732 825 2738
rect 798 2681 801 2688
rect 798 2678 806 2681
rect 798 2592 801 2628
rect 802 2548 806 2551
rect 830 2462 833 2778
rect 838 2741 841 2948
rect 886 2922 889 3178
rect 894 3002 897 3038
rect 848 2903 850 2907
rect 854 2903 857 2907
rect 862 2903 864 2907
rect 858 2868 862 2871
rect 838 2738 846 2741
rect 838 2712 841 2718
rect 848 2703 850 2707
rect 854 2703 857 2707
rect 862 2703 864 2707
rect 870 2692 873 2838
rect 894 2822 897 2998
rect 918 2961 921 2988
rect 914 2958 921 2961
rect 926 2962 929 3038
rect 942 2952 945 3138
rect 950 3122 953 3278
rect 966 3222 969 3528
rect 982 3342 985 3478
rect 974 3162 977 3168
rect 950 3002 953 3038
rect 942 2942 945 2948
rect 878 2732 881 2738
rect 850 2628 854 2631
rect 848 2503 850 2507
rect 854 2503 857 2507
rect 862 2503 864 2507
rect 838 2312 841 2468
rect 870 2362 873 2688
rect 878 2672 881 2688
rect 878 2642 881 2648
rect 886 2542 889 2788
rect 894 2782 897 2818
rect 894 2712 897 2718
rect 894 2602 897 2698
rect 878 2532 881 2538
rect 894 2382 897 2568
rect 902 2562 905 2738
rect 918 2632 921 2748
rect 910 2552 913 2558
rect 782 1862 785 1888
rect 766 1848 774 1851
rect 766 1612 769 1848
rect 790 1752 793 1898
rect 798 1762 801 2158
rect 806 1822 809 2308
rect 848 2303 850 2307
rect 854 2303 857 2307
rect 862 2303 864 2307
rect 870 2302 873 2318
rect 894 2261 897 2348
rect 890 2258 897 2261
rect 814 1742 817 1748
rect 774 1722 777 1728
rect 782 1432 785 1708
rect 798 1462 801 1658
rect 806 1532 809 1738
rect 822 1552 825 2258
rect 830 1672 833 2188
rect 848 2103 850 2107
rect 854 2103 857 2107
rect 862 2103 864 2107
rect 838 1912 841 1948
rect 848 1903 850 1907
rect 854 1903 857 1907
rect 862 1903 864 1907
rect 848 1703 850 1707
rect 854 1703 857 1707
rect 862 1703 864 1707
rect 870 1652 873 1958
rect 878 1712 881 1798
rect 886 1662 889 1988
rect 894 1952 897 2258
rect 910 2042 913 2168
rect 918 2112 921 2628
rect 926 2352 929 2588
rect 934 2502 937 2728
rect 942 2662 945 2698
rect 950 2572 953 2988
rect 958 2582 961 2738
rect 942 2482 945 2528
rect 958 2462 961 2508
rect 934 2122 937 2448
rect 966 2402 969 3078
rect 974 2932 977 3138
rect 982 2892 985 3268
rect 998 3162 1001 3168
rect 974 2662 977 2688
rect 990 2681 993 2788
rect 1014 2772 1017 2808
rect 1010 2758 1014 2761
rect 986 2678 993 2681
rect 1014 2672 1017 2728
rect 982 2628 990 2631
rect 982 2622 985 2628
rect 1006 2622 1009 2628
rect 974 2252 977 2538
rect 982 2512 985 2618
rect 1006 2492 1009 2618
rect 982 2482 985 2488
rect 990 2462 993 2468
rect 994 2348 998 2351
rect 1014 2272 1017 2668
rect 1022 2562 1025 3298
rect 1038 2712 1041 3048
rect 1046 2842 1049 2968
rect 1034 2658 1038 2661
rect 1046 2612 1049 2838
rect 1062 2762 1065 3538
rect 1070 3422 1073 3588
rect 1114 3338 1118 3341
rect 1094 3112 1097 3248
rect 1094 2872 1097 3068
rect 1054 2572 1057 2758
rect 1070 2462 1073 2858
rect 1118 2852 1121 3028
rect 1078 2672 1081 2838
rect 1134 2792 1137 3298
rect 1126 2692 1129 2788
rect 1142 2692 1145 3508
rect 1150 2762 1153 2788
rect 1086 2682 1089 2688
rect 1098 2538 1102 2541
rect 962 2138 966 2141
rect 830 1512 833 1518
rect 838 1472 841 1628
rect 848 1503 850 1507
rect 854 1503 857 1507
rect 862 1503 864 1507
rect 654 682 657 728
rect 662 702 665 818
rect 678 762 681 1048
rect 686 882 689 1178
rect 706 1138 710 1141
rect 662 262 665 698
rect 734 332 737 818
rect 578 58 585 61
rect 726 11 729 98
rect 750 72 753 718
rect 766 92 769 158
rect 774 122 777 1248
rect 782 572 785 1388
rect 790 752 793 938
rect 806 782 809 1388
rect 830 1358 838 1361
rect 830 1332 833 1358
rect 846 1352 849 1488
rect 794 488 798 491
rect 806 482 809 488
rect 814 282 817 1328
rect 848 1303 850 1307
rect 854 1303 857 1307
rect 862 1303 864 1307
rect 870 1152 873 1648
rect 886 1342 889 1378
rect 886 1182 889 1308
rect 894 1302 897 1948
rect 918 1872 921 1938
rect 950 1921 953 2008
rect 1030 1992 1033 2458
rect 1094 2272 1097 2278
rect 1074 2248 1078 2251
rect 990 1952 993 1958
rect 998 1952 1001 1958
rect 950 1918 958 1921
rect 942 1908 950 1911
rect 906 1688 910 1691
rect 918 1612 921 1848
rect 942 1842 945 1908
rect 958 1762 961 1888
rect 942 1728 950 1731
rect 942 1722 945 1728
rect 930 1718 934 1721
rect 966 1712 969 1868
rect 1038 1731 1041 2238
rect 1046 2002 1049 2248
rect 1062 1882 1065 2248
rect 1102 2162 1105 2528
rect 1118 2281 1121 2348
rect 1114 2278 1121 2281
rect 1126 2262 1129 2538
rect 1134 2452 1137 2458
rect 1126 2162 1129 2168
rect 1134 2082 1137 2438
rect 1142 2232 1145 2538
rect 1150 2192 1153 2578
rect 1158 2162 1161 3268
rect 1166 2212 1169 3468
rect 1270 3381 1273 3588
rect 1290 3518 1294 3521
rect 1270 3378 1281 3381
rect 1182 3282 1185 3318
rect 1262 3242 1265 3358
rect 1262 3162 1265 3238
rect 1234 3048 1238 3051
rect 1174 2572 1177 3038
rect 1262 2992 1265 3158
rect 1270 2982 1273 3238
rect 1254 2972 1257 2978
rect 1222 2968 1230 2971
rect 1222 2962 1225 2968
rect 1270 2942 1273 2958
rect 1242 2938 1246 2941
rect 1182 2862 1185 2888
rect 1174 2092 1177 2538
rect 1182 2092 1185 2818
rect 1198 2652 1201 2848
rect 1206 2522 1209 2868
rect 1246 2762 1249 2938
rect 1190 2372 1193 2508
rect 1198 2452 1201 2458
rect 1198 2152 1201 2348
rect 1206 2232 1209 2488
rect 1214 2472 1217 2728
rect 1034 1728 1041 1731
rect 1030 1718 1038 1721
rect 942 1652 945 1658
rect 982 1642 985 1658
rect 830 942 833 1108
rect 848 1103 850 1107
rect 854 1103 857 1107
rect 862 1103 864 1107
rect 822 722 825 908
rect 838 762 841 1088
rect 886 1042 889 1178
rect 898 1068 902 1071
rect 848 903 850 907
rect 854 903 857 907
rect 862 903 864 907
rect 886 772 889 1038
rect 838 452 841 758
rect 848 703 850 707
rect 854 703 857 707
rect 862 703 864 707
rect 848 503 850 507
rect 854 503 857 507
rect 862 503 864 507
rect 870 472 873 608
rect 906 538 910 541
rect 926 452 929 1548
rect 934 1152 937 1398
rect 942 1362 945 1508
rect 950 1342 953 1528
rect 990 1492 993 1658
rect 998 1652 1001 1668
rect 966 1312 969 1458
rect 934 1072 937 1148
rect 946 1058 950 1061
rect 958 972 961 1278
rect 966 1102 969 1308
rect 974 1072 977 1468
rect 1014 1452 1017 1668
rect 1022 1622 1025 1718
rect 1030 1602 1033 1718
rect 1038 1672 1041 1678
rect 1038 1382 1041 1448
rect 1002 1148 1006 1151
rect 958 892 961 968
rect 974 582 977 1068
rect 994 1058 998 1061
rect 1006 882 1009 938
rect 1006 732 1009 878
rect 1014 492 1017 1328
rect 1038 1142 1041 1378
rect 1046 1142 1049 1738
rect 1058 1728 1062 1731
rect 1058 1688 1062 1691
rect 1070 1552 1073 1858
rect 1150 1832 1153 2058
rect 1086 1562 1089 1798
rect 1098 1658 1102 1661
rect 1110 1492 1113 1668
rect 1150 1582 1153 1828
rect 1054 1462 1057 1468
rect 1062 1462 1065 1468
rect 1070 1342 1073 1348
rect 1062 1312 1065 1318
rect 1078 1262 1081 1418
rect 1094 1312 1097 1488
rect 1082 1138 1086 1141
rect 1022 1092 1025 1138
rect 1094 1052 1097 1298
rect 1026 868 1030 871
rect 1046 692 1049 928
rect 1094 872 1097 1048
rect 1102 1022 1105 1118
rect 1110 1082 1113 1268
rect 1118 1212 1121 1228
rect 1086 868 1094 871
rect 848 303 850 307
rect 854 303 857 307
rect 862 303 864 307
rect 848 103 850 107
rect 854 103 857 107
rect 862 103 864 107
rect 902 81 905 418
rect 974 352 977 378
rect 938 338 942 341
rect 1022 341 1025 368
rect 1018 338 1025 341
rect 1022 272 1025 278
rect 1030 182 1033 538
rect 1070 388 1078 391
rect 1070 352 1073 388
rect 1070 132 1073 178
rect 902 78 910 81
rect 1086 12 1089 868
rect 1110 542 1113 898
rect 1118 882 1121 1078
rect 1126 862 1129 1358
rect 1134 1272 1137 1458
rect 1158 1392 1161 2018
rect 1174 2012 1177 2088
rect 1182 1842 1185 2008
rect 1198 1982 1201 2138
rect 1214 2042 1217 2438
rect 1222 2382 1225 2528
rect 1230 2512 1233 2738
rect 1238 2658 1246 2661
rect 1238 2492 1241 2658
rect 1234 2428 1238 2431
rect 1230 2332 1233 2338
rect 1238 2332 1241 2358
rect 1254 2132 1257 2628
rect 1278 2562 1281 3378
rect 1286 3232 1289 3498
rect 1302 3382 1305 3528
rect 1318 3372 1321 3408
rect 1294 3262 1297 3268
rect 1286 2952 1289 2958
rect 1294 2872 1297 3248
rect 1302 2932 1305 3248
rect 1310 3242 1313 3368
rect 1318 3192 1321 3328
rect 1326 2982 1329 3288
rect 1322 2958 1326 2961
rect 1302 2922 1305 2928
rect 1302 2862 1305 2868
rect 1334 2772 1337 3588
rect 1360 3403 1362 3407
rect 1366 3403 1369 3407
rect 1374 3403 1376 3407
rect 1354 3338 1358 3341
rect 1350 3182 1353 3338
rect 1382 3322 1385 3408
rect 1360 3203 1362 3207
rect 1366 3203 1369 3207
rect 1374 3203 1376 3207
rect 1360 3003 1362 3007
rect 1366 3003 1369 3007
rect 1374 3003 1376 3007
rect 1390 3002 1393 3538
rect 1398 3322 1401 3578
rect 1418 3468 1422 3471
rect 1402 3258 1406 3261
rect 1406 3102 1409 3238
rect 1350 2812 1353 2848
rect 1360 2803 1362 2807
rect 1366 2803 1369 2807
rect 1374 2803 1376 2807
rect 1398 2762 1401 3068
rect 1406 3032 1409 3068
rect 1286 2532 1289 2618
rect 1294 2342 1297 2348
rect 1262 1992 1265 2328
rect 1270 2112 1273 2148
rect 1182 1672 1185 1808
rect 1182 1562 1185 1628
rect 1190 1532 1193 1868
rect 1134 962 1137 1198
rect 1134 862 1137 958
rect 1142 872 1145 1298
rect 1150 1252 1153 1268
rect 1158 1082 1161 1388
rect 1166 1222 1169 1488
rect 1174 1382 1177 1508
rect 1190 1491 1193 1528
rect 1186 1488 1193 1491
rect 1198 1252 1201 1878
rect 1214 1741 1217 1968
rect 1278 1952 1281 2078
rect 1294 1972 1297 2258
rect 1310 2232 1313 2278
rect 1310 2112 1313 2138
rect 1334 1992 1337 2408
rect 1342 2182 1345 2738
rect 1360 2603 1362 2607
rect 1366 2603 1369 2607
rect 1374 2603 1376 2607
rect 1360 2403 1362 2407
rect 1366 2403 1369 2407
rect 1374 2403 1376 2407
rect 1382 2352 1385 2548
rect 1354 2258 1358 2261
rect 1360 2203 1362 2207
rect 1366 2203 1369 2207
rect 1374 2203 1376 2207
rect 1360 2003 1362 2007
rect 1366 2003 1369 2007
rect 1374 2003 1376 2007
rect 1214 1738 1222 1741
rect 1206 1532 1209 1638
rect 1230 1601 1233 1688
rect 1238 1682 1241 1858
rect 1278 1792 1281 1948
rect 1302 1862 1305 1878
rect 1238 1672 1241 1678
rect 1230 1598 1238 1601
rect 1158 1042 1161 1078
rect 1154 1028 1158 1031
rect 1106 368 1110 371
rect 1110 332 1113 348
rect 1094 292 1097 328
rect 1102 252 1105 268
rect 1118 72 1121 708
rect 1142 572 1145 868
rect 1150 732 1153 838
rect 1166 782 1169 1138
rect 1198 1132 1201 1248
rect 1206 922 1209 1458
rect 1242 1328 1246 1331
rect 1246 1132 1249 1328
rect 1254 1142 1257 1608
rect 1278 1442 1281 1508
rect 1270 1342 1273 1348
rect 1262 1292 1265 1338
rect 1286 1272 1289 1588
rect 1302 1392 1305 1618
rect 1310 1482 1313 1958
rect 1310 1342 1313 1478
rect 1318 1462 1321 1988
rect 1382 1952 1385 2258
rect 1390 2172 1393 2568
rect 1390 2052 1393 2168
rect 1334 1742 1337 1868
rect 1360 1803 1362 1807
rect 1366 1803 1369 1807
rect 1374 1803 1376 1807
rect 1374 1742 1377 1758
rect 1382 1752 1385 1948
rect 1326 1622 1329 1648
rect 1334 1642 1337 1738
rect 1350 1662 1353 1668
rect 1382 1662 1385 1748
rect 1326 1482 1329 1518
rect 1270 1248 1278 1251
rect 1270 1192 1273 1248
rect 1246 1112 1249 1118
rect 1222 1081 1225 1088
rect 1218 1078 1225 1081
rect 1234 1078 1238 1081
rect 1254 1002 1257 1138
rect 1262 1122 1265 1128
rect 1270 1112 1273 1188
rect 1318 1152 1321 1458
rect 1326 1172 1329 1478
rect 1342 1302 1345 1658
rect 1360 1603 1362 1607
rect 1366 1603 1369 1607
rect 1374 1603 1376 1607
rect 1350 1492 1353 1598
rect 1382 1412 1385 1418
rect 1360 1403 1362 1407
rect 1366 1403 1369 1407
rect 1374 1403 1376 1407
rect 1350 1182 1353 1398
rect 1360 1203 1362 1207
rect 1366 1203 1369 1207
rect 1374 1203 1376 1207
rect 1318 1082 1321 1148
rect 1382 1122 1385 1198
rect 1398 1182 1401 2468
rect 1406 1552 1409 2928
rect 1414 2142 1417 3288
rect 1422 3062 1425 3118
rect 1430 3022 1433 3348
rect 1438 2938 1446 2941
rect 1422 2242 1425 2768
rect 1438 2752 1441 2938
rect 1438 2462 1441 2728
rect 1430 1892 1433 2348
rect 1438 2062 1441 2458
rect 1446 2272 1449 2278
rect 1446 2122 1449 2178
rect 1454 2122 1457 2738
rect 1430 1862 1433 1888
rect 1454 1652 1457 2118
rect 1462 2062 1465 2498
rect 1470 2472 1473 3108
rect 1478 2962 1481 3598
rect 1510 3292 1513 3598
rect 1790 3588 1798 3591
rect 1574 3402 1577 3588
rect 1478 2882 1481 2888
rect 1478 2692 1481 2868
rect 1486 2802 1489 3068
rect 1510 2922 1513 2938
rect 1518 2912 1521 3008
rect 1526 2942 1529 3158
rect 1542 2942 1545 3118
rect 1550 3062 1553 3138
rect 1550 2972 1553 2978
rect 1502 2882 1505 2888
rect 1494 2702 1497 2868
rect 1558 2862 1561 3368
rect 1478 2402 1481 2538
rect 1470 2152 1473 2398
rect 1482 2338 1486 2341
rect 1494 2271 1497 2698
rect 1518 2492 1521 2568
rect 1510 2462 1513 2488
rect 1490 2268 1497 2271
rect 1502 2272 1505 2278
rect 1470 1902 1473 1948
rect 1478 1671 1481 1688
rect 1478 1668 1486 1671
rect 1502 1671 1505 2178
rect 1510 2172 1513 2248
rect 1526 2242 1529 2778
rect 1518 2132 1521 2188
rect 1510 1872 1513 1878
rect 1518 1872 1521 2128
rect 1526 1902 1529 2078
rect 1534 1952 1537 2458
rect 1542 2432 1545 2508
rect 1550 2282 1553 2518
rect 1566 2512 1569 2988
rect 1558 2222 1561 2468
rect 1566 2442 1569 2458
rect 1558 2172 1561 2218
rect 1518 1682 1521 1868
rect 1550 1812 1553 2148
rect 1566 2022 1569 2428
rect 1566 1902 1569 1938
rect 1574 1822 1577 2828
rect 1582 2622 1585 3538
rect 1606 3422 1609 3588
rect 1598 3052 1601 3058
rect 1606 2972 1609 3418
rect 1650 3368 1654 3371
rect 1650 3268 1654 3271
rect 1614 2942 1617 3108
rect 1622 3012 1625 3038
rect 1654 2962 1657 3078
rect 1662 2982 1665 3538
rect 1750 3402 1753 3448
rect 1750 3232 1753 3398
rect 1678 3072 1681 3108
rect 1710 3102 1713 3198
rect 1734 3118 1742 3121
rect 1734 3092 1737 3118
rect 1670 2992 1673 3048
rect 1678 3042 1681 3048
rect 1686 2972 1689 3068
rect 1594 2938 1598 2941
rect 1626 2928 1630 2931
rect 1590 2722 1593 2728
rect 1590 2672 1593 2718
rect 1606 2622 1609 2848
rect 1618 2758 1622 2761
rect 1630 2552 1633 2558
rect 1582 2062 1585 2258
rect 1590 2092 1593 2378
rect 1602 2358 1606 2361
rect 1606 2152 1609 2268
rect 1606 1952 1609 2148
rect 1614 2142 1617 2148
rect 1582 1912 1585 1928
rect 1590 1892 1593 1908
rect 1598 1892 1601 1898
rect 1574 1802 1577 1818
rect 1574 1742 1577 1768
rect 1582 1742 1585 1828
rect 1590 1782 1593 1838
rect 1606 1752 1609 1948
rect 1614 1941 1617 2098
rect 1622 2082 1625 2528
rect 1638 2502 1641 2848
rect 1646 2722 1649 2728
rect 1614 1938 1622 1941
rect 1630 1938 1638 1941
rect 1630 1932 1633 1938
rect 1654 1842 1657 2958
rect 1662 2922 1665 2958
rect 1662 2692 1665 2738
rect 1670 2732 1673 2798
rect 1662 2532 1665 2608
rect 1678 2501 1681 2898
rect 1686 2742 1689 2968
rect 1726 2952 1729 2958
rect 1694 2612 1697 2898
rect 1702 2872 1705 2918
rect 1702 2752 1705 2758
rect 1702 2672 1705 2708
rect 1674 2498 1681 2501
rect 1670 2212 1673 2358
rect 1654 1742 1657 1838
rect 1642 1738 1646 1741
rect 1502 1668 1510 1671
rect 1450 1578 1457 1581
rect 1446 1452 1449 1518
rect 1454 1502 1457 1578
rect 1454 1362 1457 1368
rect 1434 1348 1438 1351
rect 1466 1348 1470 1351
rect 1406 1332 1409 1338
rect 1346 1068 1350 1071
rect 1354 1048 1358 1051
rect 1286 882 1289 1018
rect 1150 682 1153 728
rect 1142 192 1145 348
rect 1158 292 1161 438
rect 1230 392 1233 438
rect 1186 238 1190 241
rect 1194 158 1198 161
rect 1214 22 1217 148
rect 1238 142 1241 648
rect 1246 572 1249 658
rect 1278 632 1281 868
rect 1310 822 1313 878
rect 1318 872 1321 888
rect 1350 862 1353 1028
rect 1360 1003 1362 1007
rect 1366 1003 1369 1007
rect 1374 1003 1376 1007
rect 1398 832 1401 1178
rect 1406 1132 1409 1228
rect 1438 1131 1441 1148
rect 1434 1128 1441 1131
rect 1422 1052 1425 1128
rect 1438 1092 1441 1128
rect 1462 1072 1465 1218
rect 1474 1118 1478 1121
rect 1410 1048 1414 1051
rect 1422 1012 1425 1038
rect 1486 952 1489 1578
rect 1494 1392 1497 1658
rect 1554 1458 1558 1461
rect 1530 1128 1534 1131
rect 1506 1058 1510 1061
rect 1246 532 1249 568
rect 1250 458 1254 461
rect 1262 282 1265 418
rect 1278 22 1281 508
rect 1286 462 1289 468
rect 1294 282 1297 818
rect 1360 803 1362 807
rect 1366 803 1369 807
rect 1374 803 1376 807
rect 1286 162 1289 168
rect 1310 92 1313 758
rect 1360 603 1362 607
rect 1366 603 1369 607
rect 1374 603 1376 607
rect 1322 548 1326 551
rect 1366 542 1369 568
rect 1382 502 1385 788
rect 1390 552 1393 588
rect 1360 403 1362 407
rect 1366 403 1369 407
rect 1374 403 1376 407
rect 1350 382 1353 398
rect 1382 272 1385 458
rect 1390 342 1393 468
rect 1342 32 1345 208
rect 1350 202 1353 218
rect 1360 203 1362 207
rect 1366 203 1369 207
rect 1374 203 1376 207
rect 1398 162 1401 828
rect 1406 572 1409 798
rect 1414 671 1417 848
rect 1414 668 1422 671
rect 1454 652 1457 878
rect 1486 842 1489 868
rect 1494 682 1497 1038
rect 1502 872 1505 878
rect 1510 772 1513 1058
rect 1510 752 1513 758
rect 1454 602 1457 648
rect 1406 412 1409 568
rect 1430 462 1433 518
rect 1438 512 1441 548
rect 1446 502 1449 538
rect 1438 461 1441 498
rect 1438 458 1446 461
rect 1438 232 1441 238
rect 1462 132 1465 678
rect 1486 462 1489 578
rect 1510 472 1513 718
rect 1486 442 1489 458
rect 1518 452 1521 1128
rect 1526 1022 1529 1058
rect 1542 942 1545 1128
rect 1550 1002 1553 1448
rect 1558 1152 1561 1308
rect 1590 1132 1593 1668
rect 1614 1602 1617 1618
rect 1610 1548 1614 1551
rect 1622 1402 1625 1728
rect 1630 1708 1638 1711
rect 1630 1592 1633 1708
rect 1638 1632 1641 1678
rect 1630 1442 1633 1448
rect 1610 1378 1614 1381
rect 1618 1328 1625 1331
rect 1622 1312 1625 1328
rect 1622 1192 1625 1308
rect 1590 1118 1598 1121
rect 1550 952 1553 998
rect 1558 882 1561 1068
rect 1566 942 1569 1088
rect 1590 1001 1593 1118
rect 1586 998 1593 1001
rect 1590 942 1593 998
rect 1598 958 1606 961
rect 1570 848 1574 851
rect 1574 762 1577 768
rect 1542 742 1545 758
rect 1562 748 1566 751
rect 1534 582 1537 598
rect 1590 552 1593 898
rect 1598 762 1601 958
rect 1598 672 1601 688
rect 1602 668 1606 671
rect 1502 282 1505 288
rect 1518 281 1521 288
rect 1514 278 1521 281
rect 1534 272 1537 478
rect 1542 442 1545 548
rect 1550 532 1553 538
rect 1578 518 1585 521
rect 1558 462 1561 508
rect 1582 402 1585 518
rect 1590 492 1593 518
rect 1598 452 1601 588
rect 1614 552 1617 1108
rect 1622 962 1625 1188
rect 1630 812 1633 1438
rect 1646 1252 1649 1608
rect 1638 1072 1641 1118
rect 1646 1072 1649 1138
rect 1654 1052 1657 1608
rect 1662 1602 1665 1878
rect 1670 1782 1673 1868
rect 1678 1802 1681 2498
rect 1686 2182 1689 2348
rect 1686 1942 1689 1948
rect 1670 1662 1673 1778
rect 1662 1262 1665 1268
rect 1670 1112 1673 1658
rect 1678 1362 1681 1418
rect 1686 1152 1689 1848
rect 1694 1732 1697 2538
rect 1702 2182 1705 2358
rect 1710 1962 1713 2778
rect 1742 2772 1745 2808
rect 1734 2762 1737 2768
rect 1738 2748 1742 2751
rect 1742 2732 1745 2738
rect 1718 2382 1721 2708
rect 1726 2542 1729 2648
rect 1734 2542 1737 2718
rect 1750 2681 1753 3228
rect 1758 3122 1761 3588
rect 1782 3282 1785 3288
rect 1790 3172 1793 3588
rect 1802 3538 1806 3541
rect 1798 3212 1801 3398
rect 1798 3162 1801 3168
rect 1742 2678 1753 2681
rect 1718 2322 1721 2328
rect 1734 2282 1737 2288
rect 1734 2192 1737 2208
rect 1718 1962 1721 2178
rect 1734 2052 1737 2068
rect 1702 1372 1705 1888
rect 1726 1882 1729 1928
rect 1742 1892 1745 2678
rect 1758 2661 1761 2838
rect 1766 2812 1769 2818
rect 1758 2658 1766 2661
rect 1750 2262 1753 2628
rect 1758 2552 1761 2558
rect 1774 2402 1777 2558
rect 1782 2542 1785 2868
rect 1790 2812 1793 3038
rect 1798 2882 1801 3018
rect 1790 2652 1793 2788
rect 1806 2751 1809 3268
rect 1846 3022 1849 3338
rect 1862 3312 1865 3558
rect 1880 3503 1882 3507
rect 1886 3503 1889 3507
rect 1894 3503 1896 3507
rect 1874 3478 1878 3481
rect 1846 2932 1849 2938
rect 1834 2928 1841 2931
rect 1838 2922 1841 2928
rect 1798 2748 1809 2751
rect 1782 2492 1785 2508
rect 1774 2358 1782 2361
rect 1750 2122 1753 2248
rect 1766 2212 1769 2238
rect 1766 1782 1769 2178
rect 1774 2032 1777 2358
rect 1786 2268 1790 2271
rect 1782 2062 1785 2098
rect 1798 2062 1801 2748
rect 1814 2742 1817 2748
rect 1806 2728 1814 2731
rect 1806 2662 1809 2728
rect 1854 2722 1857 3148
rect 1870 3102 1873 3418
rect 1880 3303 1882 3307
rect 1886 3303 1889 3307
rect 1894 3303 1896 3307
rect 1902 3261 1905 3588
rect 1922 3348 1926 3351
rect 1898 3258 1905 3261
rect 1894 3252 1897 3258
rect 1926 3198 1934 3201
rect 1880 3103 1882 3107
rect 1886 3103 1889 3107
rect 1894 3103 1896 3107
rect 1878 2922 1881 2998
rect 1862 2832 1865 2918
rect 1902 2912 1905 2918
rect 1870 2882 1873 2908
rect 1880 2903 1882 2907
rect 1886 2903 1889 2907
rect 1894 2903 1896 2907
rect 1822 2662 1825 2678
rect 1830 2662 1833 2698
rect 1830 2552 1833 2558
rect 1818 2548 1822 2551
rect 1790 2058 1798 2061
rect 1774 1922 1777 1938
rect 1790 1822 1793 2058
rect 1798 2042 1801 2048
rect 1718 1432 1721 1518
rect 1702 1332 1705 1368
rect 1698 1268 1705 1271
rect 1702 1182 1705 1268
rect 1718 1262 1721 1328
rect 1726 1272 1729 1668
rect 1742 1512 1745 1548
rect 1730 1178 1734 1181
rect 1678 1082 1681 1148
rect 1662 1072 1665 1078
rect 1662 1052 1665 1058
rect 1638 902 1641 1038
rect 1646 772 1649 1008
rect 1654 662 1657 1048
rect 1666 998 1670 1001
rect 1718 962 1721 1018
rect 1726 962 1729 1168
rect 1726 952 1729 958
rect 1702 928 1710 931
rect 1702 812 1705 928
rect 1726 832 1729 918
rect 1710 632 1713 728
rect 1742 682 1745 1218
rect 1750 752 1753 1648
rect 1766 1202 1769 1778
rect 1790 1762 1793 1818
rect 1798 1782 1801 2038
rect 1806 2022 1809 2548
rect 1814 2332 1817 2408
rect 1814 2222 1817 2278
rect 1814 2172 1817 2218
rect 1822 2112 1825 2518
rect 1830 2032 1833 2478
rect 1838 2452 1841 2668
rect 1850 2538 1854 2541
rect 1862 2522 1865 2828
rect 1870 2752 1873 2758
rect 1880 2703 1882 2707
rect 1886 2703 1889 2707
rect 1894 2703 1896 2707
rect 1870 2692 1873 2698
rect 1890 2608 1894 2611
rect 1880 2503 1882 2507
rect 1886 2503 1889 2507
rect 1894 2503 1896 2507
rect 1838 2372 1841 2448
rect 1838 2251 1841 2348
rect 1854 2342 1857 2348
rect 1862 2308 1870 2311
rect 1846 2272 1849 2308
rect 1854 2252 1857 2288
rect 1862 2272 1865 2308
rect 1880 2303 1882 2307
rect 1886 2303 1889 2307
rect 1894 2303 1896 2307
rect 1838 2248 1846 2251
rect 1902 2182 1905 2858
rect 1910 2562 1913 3158
rect 1926 3072 1929 3198
rect 1926 2642 1929 3028
rect 1910 2502 1913 2558
rect 1914 2488 1918 2491
rect 1926 2452 1929 2638
rect 1934 2632 1937 3138
rect 1958 2972 1961 3598
rect 2074 3588 2081 3591
rect 2002 3538 2006 3541
rect 1974 3522 1977 3528
rect 1942 2712 1945 2948
rect 1830 1952 1833 2028
rect 1838 2012 1841 2018
rect 1846 1952 1849 2178
rect 1854 2152 1857 2158
rect 1926 2152 1929 2158
rect 1862 2052 1865 2108
rect 1870 2071 1873 2118
rect 1880 2103 1882 2107
rect 1886 2103 1889 2107
rect 1894 2103 1896 2107
rect 1910 2082 1913 2138
rect 1870 2068 1878 2071
rect 1926 2062 1929 2088
rect 1934 2062 1937 2548
rect 1942 2462 1945 2708
rect 1958 2682 1961 2728
rect 1950 2462 1953 2578
rect 1958 2472 1961 2628
rect 1806 1902 1809 1918
rect 1774 1662 1777 1688
rect 1782 1642 1785 1668
rect 1806 1662 1809 1758
rect 1846 1612 1849 1948
rect 1862 1582 1865 2048
rect 1926 1982 1929 2058
rect 1942 2052 1945 2308
rect 1880 1903 1882 1907
rect 1886 1903 1889 1907
rect 1894 1903 1896 1907
rect 1870 1702 1873 1728
rect 1880 1703 1882 1707
rect 1886 1703 1889 1707
rect 1894 1703 1896 1707
rect 1902 1702 1905 1728
rect 1910 1712 1913 1768
rect 1790 1402 1793 1538
rect 1798 1462 1801 1538
rect 1870 1532 1873 1698
rect 1910 1682 1913 1688
rect 1918 1672 1921 1718
rect 1926 1612 1929 1718
rect 1880 1503 1882 1507
rect 1886 1503 1889 1507
rect 1894 1503 1896 1507
rect 1902 1482 1905 1558
rect 1942 1492 1945 2048
rect 1950 1912 1953 2458
rect 1958 2352 1961 2468
rect 1966 2392 1969 3128
rect 1974 2972 1977 2978
rect 1982 2782 1985 3528
rect 2022 3312 2025 3468
rect 1998 3052 2001 3058
rect 2006 3052 2009 3078
rect 1990 2762 1993 2768
rect 1990 2752 1993 2758
rect 1958 2092 1961 2218
rect 1966 2122 1969 2158
rect 1974 2062 1977 2208
rect 1982 2172 1985 2718
rect 1990 2262 1993 2678
rect 1998 2092 2001 3018
rect 2014 2982 2017 3298
rect 2022 3072 2025 3148
rect 2010 2968 2017 2971
rect 2006 2932 2009 2938
rect 2014 2932 2017 2968
rect 2022 2872 2025 3068
rect 2030 2982 2033 3088
rect 2038 3082 2041 3128
rect 2062 3052 2065 3198
rect 2050 2978 2054 2981
rect 2014 2752 2017 2868
rect 2022 2742 2025 2868
rect 2030 2742 2033 2748
rect 2030 2322 2033 2358
rect 2030 2312 2033 2318
rect 2006 2272 2009 2298
rect 2006 2252 2009 2268
rect 2014 2221 2017 2228
rect 2010 2218 2017 2221
rect 2022 2212 2025 2228
rect 2022 2172 2025 2188
rect 1974 1942 1977 2058
rect 1998 1952 2001 2088
rect 1958 1841 1961 1848
rect 1954 1838 1961 1841
rect 1946 1488 1950 1491
rect 1878 1452 1881 1478
rect 1910 1462 1913 1478
rect 1910 1452 1913 1458
rect 1942 1442 1945 1448
rect 1886 1392 1889 1408
rect 1882 1358 1886 1361
rect 1774 1182 1777 1358
rect 1838 1302 1841 1318
rect 1834 1298 1838 1301
rect 1766 1082 1769 1148
rect 1774 1052 1777 1158
rect 1766 1022 1769 1028
rect 1766 882 1769 1018
rect 1766 762 1769 878
rect 1774 872 1777 1048
rect 1646 562 1649 588
rect 1606 482 1609 488
rect 1546 338 1550 341
rect 1522 268 1526 271
rect 1534 262 1537 268
rect 1530 248 1534 251
rect 1558 242 1561 298
rect 1614 272 1617 528
rect 1718 502 1721 578
rect 1726 502 1729 648
rect 1750 472 1753 748
rect 1790 532 1793 548
rect 1578 268 1582 271
rect 1590 182 1593 268
rect 1622 252 1625 288
rect 1614 182 1617 248
rect 1622 202 1625 218
rect 1646 92 1649 218
rect 1654 172 1657 178
rect 1662 72 1665 178
rect 1686 152 1689 358
rect 1702 251 1705 268
rect 1702 248 1710 251
rect 1742 142 1745 328
rect 1750 272 1753 468
rect 1766 252 1769 418
rect 1774 251 1777 288
rect 1774 248 1782 251
rect 1790 102 1793 528
rect 1798 482 1801 908
rect 1806 762 1809 1178
rect 1814 1142 1817 1178
rect 1846 1082 1849 1268
rect 1870 1162 1873 1358
rect 1880 1303 1882 1307
rect 1886 1303 1889 1307
rect 1894 1303 1896 1307
rect 1834 1028 1838 1031
rect 1814 942 1817 988
rect 1826 948 1830 951
rect 1846 942 1849 1078
rect 1854 972 1857 1118
rect 1870 1012 1873 1108
rect 1880 1103 1882 1107
rect 1886 1103 1889 1107
rect 1894 1103 1896 1107
rect 1902 1082 1905 1278
rect 1850 938 1854 941
rect 1826 848 1830 851
rect 1814 822 1817 848
rect 1806 82 1809 678
rect 1814 472 1817 738
rect 1826 468 1830 471
rect 1814 412 1817 468
rect 1838 362 1841 618
rect 1846 482 1849 898
rect 1870 862 1873 948
rect 1880 903 1882 907
rect 1886 903 1889 907
rect 1894 903 1896 907
rect 1894 882 1897 888
rect 1858 798 1862 801
rect 1854 492 1857 778
rect 1862 692 1865 798
rect 1870 772 1873 798
rect 1880 703 1882 707
rect 1886 703 1889 707
rect 1894 703 1896 707
rect 1880 503 1882 507
rect 1886 503 1889 507
rect 1894 503 1896 507
rect 1902 492 1905 1078
rect 1910 952 1913 1318
rect 1934 1191 1937 1308
rect 1946 1268 1950 1271
rect 1930 1188 1937 1191
rect 1922 948 1929 951
rect 1910 702 1913 878
rect 1926 852 1929 948
rect 1934 832 1937 1068
rect 1950 832 1953 1128
rect 1958 1082 1961 1558
rect 1966 1492 1969 1908
rect 2006 1792 2009 2038
rect 2030 1932 2033 2298
rect 2030 1882 2033 1928
rect 1970 1188 1974 1191
rect 1966 972 1969 1138
rect 1958 962 1961 968
rect 1958 892 1961 918
rect 1966 862 1969 968
rect 1974 942 1977 958
rect 1918 712 1921 738
rect 1926 662 1929 668
rect 1862 352 1865 478
rect 1934 472 1937 738
rect 1942 632 1945 828
rect 1950 672 1953 738
rect 1974 681 1977 868
rect 1982 842 1985 1738
rect 1990 1722 1993 1728
rect 2038 1592 2041 2718
rect 2046 2512 2049 2898
rect 2054 2882 2057 2968
rect 2062 2942 2065 3048
rect 2070 2982 2073 3568
rect 2078 3162 2081 3588
rect 2126 3462 2129 3558
rect 2166 3342 2169 3538
rect 2218 3418 2222 3421
rect 2070 2872 2073 2938
rect 2078 2862 2081 3058
rect 2102 2982 2105 3038
rect 2110 3032 2113 3338
rect 2118 3042 2121 3118
rect 2126 3102 2129 3318
rect 2166 3242 2169 3338
rect 2126 3002 2129 3088
rect 2134 2982 2137 3058
rect 2118 2912 2121 2978
rect 2130 2938 2134 2941
rect 2134 2928 2142 2931
rect 2134 2912 2137 2928
rect 2066 2858 2070 2861
rect 2078 2692 2081 2858
rect 2094 2812 2097 2878
rect 2142 2812 2145 2858
rect 2150 2822 2153 3158
rect 2162 3058 2169 3061
rect 2166 3052 2169 3058
rect 2190 2972 2193 3228
rect 2198 3132 2201 3328
rect 2230 3162 2233 3588
rect 2394 3538 2398 3541
rect 2238 3512 2241 3518
rect 2270 3512 2273 3528
rect 2266 3458 2270 3461
rect 2278 3392 2281 3528
rect 2306 3328 2313 3331
rect 2298 3318 2302 3321
rect 2226 3158 2230 3161
rect 2198 2892 2201 3128
rect 2226 3108 2230 3111
rect 2238 3052 2241 3128
rect 2246 3102 2249 3318
rect 2310 3202 2313 3328
rect 2238 2992 2241 3048
rect 2218 2968 2222 2971
rect 2206 2922 2209 2928
rect 2162 2858 2166 2861
rect 2046 1692 2049 2288
rect 2054 1562 2057 1928
rect 2062 1692 2065 2558
rect 2078 2522 2081 2688
rect 2110 2662 2113 2708
rect 2118 2672 2121 2788
rect 2142 2712 2145 2808
rect 2070 1762 2073 1798
rect 1998 1242 2001 1308
rect 1990 1032 1993 1038
rect 1998 781 2001 1238
rect 1970 678 1977 681
rect 1990 778 2001 781
rect 1950 542 1953 668
rect 1958 662 1961 668
rect 1946 468 1950 471
rect 1974 432 1977 448
rect 1842 338 1846 341
rect 1870 312 1873 378
rect 1942 352 1945 368
rect 1880 303 1882 307
rect 1886 303 1889 307
rect 1894 303 1896 307
rect 1910 272 1913 288
rect 1934 282 1937 288
rect 1950 262 1953 348
rect 1962 258 1966 261
rect 1842 238 1846 241
rect 1880 103 1882 107
rect 1886 103 1889 107
rect 1894 103 1896 107
rect 1926 22 1929 248
rect 1950 242 1953 258
rect 1974 252 1977 338
rect 1990 182 1993 778
rect 1998 652 2001 728
rect 2022 682 2025 1528
rect 2038 1222 2041 1458
rect 2058 1448 2062 1451
rect 2078 1362 2081 1438
rect 2062 1332 2065 1348
rect 2086 1292 2089 2248
rect 2094 2152 2097 2158
rect 2094 2132 2097 2148
rect 2102 1882 2105 2418
rect 2118 2282 2121 2548
rect 2126 1932 2129 2618
rect 2142 2312 2145 2708
rect 2154 2668 2158 2671
rect 2150 2532 2153 2658
rect 2150 2452 2153 2498
rect 2150 2262 2153 2328
rect 2158 2252 2161 2598
rect 2166 2542 2169 2778
rect 2206 2612 2209 2708
rect 2214 2642 2217 2858
rect 2222 2822 2225 2858
rect 2150 2182 2153 2198
rect 2166 2071 2169 2368
rect 2178 2268 2182 2271
rect 2174 2192 2177 2228
rect 2206 2142 2209 2448
rect 2214 2262 2217 2638
rect 2222 2202 2225 2818
rect 2246 2742 2249 3098
rect 2254 3072 2257 3148
rect 2294 3142 2297 3148
rect 2306 3138 2310 3141
rect 2254 2812 2257 3038
rect 2262 2882 2265 3058
rect 2270 3042 2273 3058
rect 2278 3032 2281 3088
rect 2286 3082 2289 3098
rect 2270 2922 2273 2948
rect 2278 2862 2281 3028
rect 2286 2882 2289 3078
rect 2246 2582 2249 2688
rect 2254 2672 2257 2788
rect 2270 2682 2273 2688
rect 2278 2652 2281 2858
rect 2278 2612 2281 2648
rect 2242 2528 2246 2531
rect 2206 2122 2209 2138
rect 2162 2068 2169 2071
rect 2182 2072 2185 2078
rect 2182 2052 2185 2068
rect 2206 2052 2209 2098
rect 2214 2052 2217 2118
rect 2146 2048 2153 2051
rect 2150 1992 2153 2048
rect 2126 1922 2129 1928
rect 2094 1878 2102 1881
rect 2094 1672 2097 1878
rect 2118 1772 2121 1908
rect 2174 1872 2177 1888
rect 2198 1872 2201 1878
rect 2126 1542 2129 1718
rect 2134 1702 2137 1728
rect 2166 1362 2169 1388
rect 2094 1352 2097 1358
rect 2126 1328 2134 1331
rect 2126 1292 2129 1328
rect 2150 1172 2153 1328
rect 2030 1142 2033 1148
rect 2038 1118 2046 1121
rect 2114 1118 2118 1121
rect 2038 1112 2041 1118
rect 2054 1082 2057 1098
rect 2086 1082 2089 1088
rect 2118 1052 2121 1118
rect 2126 1092 2129 1108
rect 2058 938 2062 941
rect 2062 912 2065 928
rect 2058 868 2062 871
rect 2034 848 2041 851
rect 2038 842 2041 848
rect 2010 648 2017 651
rect 2014 612 2017 648
rect 2014 462 2017 608
rect 2014 362 2017 368
rect 2022 332 2025 608
rect 2038 572 2041 658
rect 2062 642 2065 758
rect 2062 591 2065 638
rect 2062 588 2070 591
rect 2078 552 2081 908
rect 2102 822 2105 1048
rect 2142 1002 2145 1158
rect 2150 991 2153 1148
rect 2166 1112 2169 1158
rect 2174 1122 2177 1488
rect 2182 1072 2185 1078
rect 2190 1062 2193 1348
rect 2206 1082 2209 1958
rect 2222 1402 2225 2198
rect 2230 2162 2233 2208
rect 2230 2002 2233 2068
rect 2230 1572 2233 1678
rect 2238 1332 2241 2528
rect 2246 2202 2249 2408
rect 2258 2278 2262 2281
rect 2278 2242 2281 2608
rect 2286 2042 2289 2758
rect 2294 2642 2297 3038
rect 2302 2862 2305 3058
rect 2318 2992 2321 3348
rect 2326 3132 2329 3138
rect 2310 2922 2313 2968
rect 2318 2912 2321 2938
rect 2294 2532 2297 2588
rect 2310 2442 2313 2848
rect 2294 2172 2297 2258
rect 2302 2071 2305 2428
rect 2314 2338 2318 2341
rect 2310 2082 2313 2268
rect 2302 2068 2313 2071
rect 2310 2062 2313 2068
rect 2262 1842 2265 1958
rect 2286 1892 2289 2038
rect 2310 1942 2313 2058
rect 2318 1992 2321 2008
rect 2274 1878 2278 1881
rect 2262 1352 2265 1838
rect 2274 1778 2278 1781
rect 2294 1742 2297 1898
rect 2302 1872 2305 1878
rect 2294 1682 2297 1738
rect 2310 1452 2313 1938
rect 2326 1912 2329 3008
rect 2334 2872 2337 3438
rect 2346 2928 2350 2931
rect 2350 2872 2353 2908
rect 2358 2852 2361 3318
rect 2374 3312 2377 3408
rect 2384 3403 2386 3407
rect 2390 3403 2393 3407
rect 2398 3403 2400 3407
rect 2406 3362 2409 3588
rect 2574 3532 2577 3538
rect 2490 3528 2497 3531
rect 2494 3522 2497 3528
rect 2574 3462 2577 3468
rect 2546 3458 2550 3461
rect 2558 3432 2561 3448
rect 2384 3203 2386 3207
rect 2390 3203 2393 3207
rect 2398 3203 2400 3207
rect 2334 2842 2337 2848
rect 2350 2772 2353 2798
rect 2358 2752 2361 2848
rect 2366 2682 2369 3048
rect 2384 3003 2386 3007
rect 2390 3003 2393 3007
rect 2398 3003 2400 3007
rect 2374 2932 2377 2938
rect 2390 2862 2393 2868
rect 2384 2803 2386 2807
rect 2390 2803 2393 2807
rect 2398 2803 2400 2807
rect 2374 2752 2377 2798
rect 2398 2682 2401 2708
rect 2406 2672 2409 2718
rect 2414 2712 2417 3418
rect 2550 3262 2553 3368
rect 2666 3308 2670 3311
rect 2870 3282 2873 3508
rect 2904 3503 2906 3507
rect 2910 3503 2913 3507
rect 2918 3503 2920 3507
rect 2926 3502 2929 3518
rect 2894 3452 2897 3478
rect 2886 3358 2894 3361
rect 2442 3058 2446 3061
rect 2422 2692 2425 3048
rect 2454 2972 2457 3118
rect 2470 3112 2473 3128
rect 2462 3052 2465 3058
rect 2454 2872 2457 2968
rect 2462 2952 2465 3048
rect 2502 2932 2505 2938
rect 2470 2872 2473 2928
rect 2418 2648 2422 2651
rect 2406 2612 2409 2648
rect 2384 2603 2386 2607
rect 2390 2603 2393 2607
rect 2398 2603 2400 2607
rect 2406 2512 2409 2548
rect 2422 2502 2425 2648
rect 2438 2531 2441 2858
rect 2454 2762 2457 2868
rect 2446 2702 2449 2718
rect 2438 2528 2449 2531
rect 2334 2328 2342 2331
rect 2334 2322 2337 2328
rect 2342 1882 2345 2128
rect 2350 2052 2353 2348
rect 2358 2212 2361 2358
rect 2366 1982 2369 2498
rect 2418 2488 2422 2491
rect 2384 2403 2386 2407
rect 2390 2403 2393 2407
rect 2398 2403 2400 2407
rect 2410 2338 2414 2341
rect 2422 2331 2425 2388
rect 2438 2332 2441 2518
rect 2422 2328 2430 2331
rect 2374 2262 2377 2268
rect 2384 2203 2386 2207
rect 2390 2203 2393 2207
rect 2398 2203 2400 2207
rect 2406 2012 2409 2038
rect 2384 2003 2386 2007
rect 2390 2003 2393 2007
rect 2398 2003 2400 2007
rect 2346 1858 2350 1861
rect 2318 1782 2321 1788
rect 2270 1362 2273 1368
rect 2270 1292 2273 1358
rect 2278 1332 2281 1338
rect 2294 1282 2297 1288
rect 2214 1132 2217 1138
rect 2178 1058 2182 1061
rect 2142 988 2153 991
rect 2122 978 2126 981
rect 2122 818 2126 821
rect 2102 732 2105 818
rect 2134 792 2137 818
rect 2102 652 2105 658
rect 2086 602 2089 628
rect 2142 602 2145 988
rect 2166 981 2169 1008
rect 2162 978 2169 981
rect 2170 948 2177 951
rect 2150 782 2153 798
rect 2174 781 2177 948
rect 2182 802 2185 998
rect 2202 928 2206 931
rect 2190 902 2193 908
rect 2222 812 2225 1218
rect 2214 792 2217 808
rect 2174 778 2182 781
rect 2214 781 2217 788
rect 2214 778 2222 781
rect 2174 702 2177 778
rect 2178 658 2185 661
rect 2030 352 2033 428
rect 2046 382 2049 388
rect 2030 292 2033 348
rect 1954 168 1958 171
rect 2014 32 2017 198
rect 2038 62 2041 378
rect 2046 192 2049 338
rect 2054 282 2057 498
rect 2086 442 2089 568
rect 2094 492 2097 598
rect 2158 562 2161 568
rect 2182 552 2185 658
rect 2134 522 2137 538
rect 2182 472 2185 548
rect 2206 481 2209 608
rect 2230 562 2233 648
rect 2238 622 2241 1268
rect 2246 642 2249 1258
rect 2294 1168 2302 1171
rect 2294 1072 2297 1168
rect 2302 1112 2305 1148
rect 2254 752 2257 888
rect 2262 752 2265 848
rect 2254 692 2257 748
rect 2266 678 2270 681
rect 2254 632 2257 678
rect 2278 672 2281 948
rect 2286 942 2289 948
rect 2286 772 2289 778
rect 2294 692 2297 768
rect 2302 562 2305 768
rect 2310 652 2313 1448
rect 2326 1322 2329 1358
rect 2318 1222 2321 1248
rect 2334 1182 2337 1788
rect 2350 1652 2353 1848
rect 2358 1822 2361 1968
rect 2374 1962 2377 1998
rect 2406 1912 2409 1948
rect 2414 1942 2417 2098
rect 2422 2082 2425 2288
rect 2438 2282 2441 2328
rect 2446 2262 2449 2528
rect 2430 2162 2433 2238
rect 2446 2142 2449 2158
rect 2430 2082 2433 2088
rect 2438 2042 2441 2128
rect 2430 1892 2433 1938
rect 2446 1932 2449 2078
rect 2454 1962 2457 2708
rect 2462 2582 2465 2808
rect 2470 2742 2473 2868
rect 2462 2542 2465 2558
rect 2470 2542 2473 2738
rect 2470 2482 2473 2538
rect 2462 2222 2465 2448
rect 2478 2332 2481 2728
rect 2486 2402 2489 2908
rect 2470 2282 2473 2318
rect 2482 2268 2486 2271
rect 2478 2171 2481 2248
rect 2474 2168 2481 2171
rect 2462 1972 2465 2168
rect 2462 1942 2465 1948
rect 2370 1868 2374 1871
rect 2414 1852 2417 1858
rect 2406 1812 2409 1838
rect 2384 1803 2386 1807
rect 2390 1803 2393 1807
rect 2398 1803 2400 1807
rect 2386 1758 2390 1761
rect 2366 1742 2369 1748
rect 2374 1742 2377 1758
rect 2398 1712 2401 1718
rect 2370 1688 2374 1691
rect 2374 1652 2377 1688
rect 2384 1603 2386 1607
rect 2390 1603 2393 1607
rect 2398 1603 2400 1607
rect 2366 1452 2369 1598
rect 2384 1403 2386 1407
rect 2390 1403 2393 1407
rect 2398 1403 2400 1407
rect 2342 1272 2345 1298
rect 2350 1162 2353 1278
rect 2374 1272 2377 1338
rect 2406 1212 2409 1668
rect 2414 1462 2417 1848
rect 2430 1792 2433 1888
rect 2438 1882 2441 1888
rect 2422 1422 2425 1438
rect 2384 1203 2386 1207
rect 2390 1203 2393 1207
rect 2398 1203 2400 1207
rect 2422 1202 2425 1418
rect 2446 1282 2449 1928
rect 2454 1862 2457 1878
rect 2454 1842 2457 1848
rect 2462 1772 2465 1938
rect 2470 1452 2473 2058
rect 2478 2032 2481 2168
rect 2494 2102 2497 2708
rect 2518 2582 2521 3138
rect 2506 2558 2513 2561
rect 2510 2552 2513 2558
rect 2494 2042 2497 2048
rect 2502 1952 2505 2548
rect 2510 2522 2513 2548
rect 2526 2352 2529 3018
rect 2550 2972 2553 3258
rect 2886 3252 2889 3358
rect 2904 3303 2906 3307
rect 2910 3303 2913 3307
rect 2918 3303 2920 3307
rect 2926 3302 2929 3328
rect 2902 3242 2905 3268
rect 2590 3122 2593 3158
rect 2574 2992 2577 3078
rect 2582 3002 2585 3068
rect 2598 3042 2601 3138
rect 2610 3058 2614 3061
rect 2550 2832 2553 2848
rect 2550 2602 2553 2828
rect 2542 2482 2545 2508
rect 2546 2258 2550 2261
rect 2510 2162 2513 2168
rect 2530 2158 2534 2161
rect 2526 2062 2529 2138
rect 2542 2102 2545 2118
rect 2526 1981 2529 2058
rect 2550 1992 2553 2128
rect 2522 1978 2529 1981
rect 2478 1731 2481 1928
rect 2510 1772 2513 1978
rect 2478 1728 2486 1731
rect 2486 1662 2489 1678
rect 2486 1332 2489 1478
rect 2502 1462 2505 1528
rect 2502 1362 2505 1388
rect 2326 1082 2329 1158
rect 2374 1152 2377 1178
rect 2374 1002 2377 1038
rect 2384 1003 2386 1007
rect 2390 1003 2393 1007
rect 2398 1003 2400 1007
rect 2374 952 2377 998
rect 2342 782 2345 948
rect 2366 932 2369 948
rect 2390 932 2393 958
rect 2422 951 2425 1168
rect 2430 1152 2433 1178
rect 2438 1122 2441 1148
rect 2454 1142 2457 1328
rect 2418 948 2425 951
rect 2366 881 2369 898
rect 2366 878 2374 881
rect 2384 803 2386 807
rect 2390 803 2393 807
rect 2398 803 2400 807
rect 2382 722 2385 728
rect 2338 658 2342 661
rect 2206 478 2214 481
rect 2086 342 2089 438
rect 2062 282 2065 288
rect 2094 22 2097 378
rect 2110 281 2113 468
rect 2254 462 2257 558
rect 2318 462 2321 638
rect 2334 542 2337 558
rect 2250 458 2254 461
rect 2134 282 2137 388
rect 2110 278 2118 281
rect 2142 152 2145 378
rect 2150 142 2153 288
rect 2174 172 2177 438
rect 2190 262 2193 388
rect 2206 292 2209 388
rect 2230 302 2233 328
rect 2222 292 2225 298
rect 2206 282 2209 288
rect 2238 281 2241 418
rect 2246 362 2249 378
rect 2274 338 2278 341
rect 2234 278 2241 281
rect 2190 172 2193 238
rect 2198 182 2201 278
rect 2102 72 2105 88
rect 2206 72 2209 228
rect 2214 202 2217 278
rect 2230 151 2233 158
rect 2222 148 2233 151
rect 2222 142 2225 148
rect 2238 142 2241 248
rect 2286 202 2289 338
rect 2310 282 2313 358
rect 2326 342 2329 348
rect 2334 342 2337 448
rect 2342 422 2345 658
rect 2350 532 2353 718
rect 2406 712 2409 848
rect 2366 622 2369 648
rect 2414 642 2417 908
rect 2422 772 2425 878
rect 2430 862 2433 1068
rect 2454 1062 2457 1138
rect 2442 1048 2446 1051
rect 2462 811 2465 1178
rect 2486 1172 2489 1328
rect 2510 1322 2513 1368
rect 2518 1262 2521 1958
rect 2558 1862 2561 2768
rect 2566 1982 2569 2068
rect 2574 1962 2577 2988
rect 2582 2892 2585 2998
rect 2618 2978 2625 2981
rect 2582 2492 2585 2858
rect 2598 2582 2601 2838
rect 2606 2761 2609 2928
rect 2622 2872 2625 2978
rect 2630 2792 2633 3168
rect 2606 2758 2614 2761
rect 2590 2412 2593 2538
rect 2598 2502 2601 2528
rect 2606 2482 2609 2518
rect 2598 2192 2601 2378
rect 2614 2372 2617 2548
rect 2622 2342 2625 2478
rect 2638 2372 2641 2858
rect 2654 2852 2657 3038
rect 2662 2932 2665 3028
rect 2662 2852 2665 2858
rect 2646 2602 2649 2678
rect 2654 2462 2657 2638
rect 2606 2202 2609 2308
rect 2626 2268 2630 2271
rect 2614 2152 2617 2248
rect 2654 2152 2657 2458
rect 2662 2182 2665 2848
rect 2670 2752 2673 3178
rect 2682 3118 2686 3121
rect 2694 2882 2697 3048
rect 2706 2938 2710 2941
rect 2774 2932 2777 3128
rect 2904 3103 2906 3107
rect 2910 3103 2913 3107
rect 2918 3103 2920 3107
rect 2694 2852 2697 2868
rect 2678 2798 2686 2801
rect 2670 2162 2673 2598
rect 2678 2512 2681 2798
rect 2694 2672 2697 2698
rect 2686 2652 2689 2668
rect 2686 2162 2689 2638
rect 2702 2442 2705 2698
rect 2710 2592 2713 2858
rect 2726 2852 2729 2898
rect 2806 2882 2809 3088
rect 2822 2882 2825 2958
rect 2722 2768 2729 2771
rect 2710 2382 2713 2468
rect 2718 2272 2721 2678
rect 2726 2662 2729 2768
rect 2770 2708 2774 2711
rect 2734 2552 2737 2668
rect 2754 2638 2758 2641
rect 2590 2092 2593 2118
rect 2606 2092 2609 2128
rect 2582 2062 2585 2078
rect 2586 2058 2590 2061
rect 2598 2042 2601 2088
rect 2614 2062 2617 2148
rect 2530 1858 2534 1861
rect 2566 1832 2569 1938
rect 2526 1742 2529 1758
rect 2566 1742 2569 1828
rect 2550 1692 2553 1728
rect 2574 1652 2577 1768
rect 2598 1552 2601 1938
rect 2526 1322 2529 1548
rect 2594 1488 2598 1491
rect 2566 1262 2569 1368
rect 2478 1162 2481 1168
rect 2498 1158 2502 1161
rect 2486 1132 2489 1138
rect 2478 1128 2486 1131
rect 2470 1112 2473 1118
rect 2478 1102 2481 1128
rect 2474 1068 2478 1071
rect 2486 1062 2489 1118
rect 2518 1082 2521 1118
rect 2494 871 2497 998
rect 2502 882 2505 1078
rect 2526 952 2529 1208
rect 2534 962 2537 1248
rect 2542 941 2545 1258
rect 2574 1192 2577 1478
rect 2590 1472 2593 1478
rect 2606 1471 2609 1488
rect 2602 1468 2609 1471
rect 2554 1128 2558 1131
rect 2558 1042 2561 1058
rect 2574 1052 2577 1058
rect 2558 962 2561 1028
rect 2566 1002 2569 1048
rect 2574 1002 2577 1048
rect 2566 962 2569 998
rect 2574 972 2577 978
rect 2582 952 2585 1288
rect 2542 938 2553 941
rect 2494 868 2502 871
rect 2514 868 2518 871
rect 2534 832 2537 938
rect 2458 808 2465 811
rect 2430 752 2433 798
rect 2446 682 2449 698
rect 2374 602 2377 618
rect 2384 603 2386 607
rect 2390 603 2393 607
rect 2398 603 2400 607
rect 2366 532 2369 588
rect 2366 442 2369 458
rect 2374 442 2377 588
rect 2446 502 2449 548
rect 2382 462 2385 478
rect 2446 472 2449 478
rect 2378 438 2382 441
rect 2384 403 2386 407
rect 2390 403 2393 407
rect 2398 403 2400 407
rect 2350 342 2353 348
rect 2374 342 2377 358
rect 2398 262 2401 388
rect 2418 338 2425 341
rect 2384 203 2386 207
rect 2390 203 2393 207
rect 2398 203 2400 207
rect 2422 192 2425 338
rect 2430 172 2433 388
rect 2438 291 2441 298
rect 2438 288 2446 291
rect 2454 282 2457 528
rect 2462 452 2465 778
rect 2478 732 2481 828
rect 2486 752 2489 808
rect 2494 792 2497 798
rect 2518 752 2521 768
rect 2498 748 2502 751
rect 2486 742 2489 748
rect 2478 692 2481 728
rect 2470 672 2473 688
rect 2490 648 2494 651
rect 2462 342 2465 408
rect 2470 302 2473 478
rect 2486 462 2489 598
rect 2478 292 2481 298
rect 2470 222 2473 268
rect 2478 192 2481 218
rect 2474 188 2478 191
rect 2254 82 2257 158
rect 2486 112 2489 438
rect 2494 352 2497 478
rect 2502 432 2505 678
rect 2518 602 2521 728
rect 2518 542 2521 598
rect 2526 592 2529 618
rect 2502 92 2505 428
rect 2510 362 2513 368
rect 2526 292 2529 378
rect 2534 332 2537 598
rect 2542 402 2545 488
rect 2550 452 2553 938
rect 2582 862 2585 908
rect 2582 652 2585 758
rect 2590 552 2593 1468
rect 2614 1262 2617 1948
rect 2622 1942 2625 2088
rect 2630 1822 2633 1948
rect 2646 1852 2649 2108
rect 2670 2042 2673 2068
rect 2698 2058 2705 2061
rect 2682 2038 2686 2041
rect 2630 1752 2633 1818
rect 2646 1662 2649 1728
rect 2598 1072 2601 1118
rect 2606 1082 2609 1168
rect 2614 1122 2617 1258
rect 2602 1058 2606 1061
rect 2622 1061 2625 1238
rect 2614 1058 2625 1061
rect 2598 902 2601 968
rect 2614 902 2617 1058
rect 2630 1052 2633 1278
rect 2654 1262 2657 1858
rect 2662 1582 2665 1878
rect 2670 1742 2673 1748
rect 2678 1472 2681 1808
rect 2686 1742 2689 1888
rect 2686 1642 2689 1658
rect 2678 1312 2681 1328
rect 2678 1282 2681 1308
rect 2646 1201 2649 1218
rect 2642 1198 2649 1201
rect 2638 1062 2641 1158
rect 2662 1131 2665 1178
rect 2662 1128 2670 1131
rect 2622 1048 2630 1051
rect 2622 932 2625 1048
rect 2630 952 2633 958
rect 2646 932 2649 1078
rect 2662 992 2665 1118
rect 2670 1072 2673 1088
rect 2654 948 2662 951
rect 2634 918 2638 921
rect 2622 762 2625 868
rect 2654 852 2657 948
rect 2678 942 2681 1148
rect 2686 962 2689 1638
rect 2694 1512 2697 1968
rect 2702 1812 2705 2058
rect 2710 1952 2713 2148
rect 2710 1792 2713 1918
rect 2710 1772 2713 1788
rect 2718 1742 2721 2138
rect 2726 1942 2729 2428
rect 2734 2142 2737 2548
rect 2742 2462 2745 2628
rect 2762 2568 2766 2571
rect 2706 1738 2710 1741
rect 2718 1692 2721 1728
rect 2710 1512 2713 1688
rect 2710 1491 2713 1498
rect 2710 1488 2718 1491
rect 2726 1462 2729 1928
rect 2734 1562 2737 2088
rect 2742 2052 2745 2338
rect 2742 1682 2745 1948
rect 2750 1932 2753 2138
rect 2758 1932 2761 1948
rect 2766 1862 2769 2118
rect 2774 2062 2777 2648
rect 2790 2622 2793 2878
rect 2798 2742 2801 2768
rect 2790 2572 2793 2578
rect 2798 2572 2801 2738
rect 2782 2432 2785 2568
rect 2798 2562 2801 2568
rect 2814 2522 2817 2718
rect 2822 2641 2825 2688
rect 2830 2652 2833 2878
rect 2862 2722 2865 2808
rect 2838 2642 2841 2668
rect 2822 2638 2830 2641
rect 2806 2332 2809 2338
rect 2790 2152 2793 2328
rect 2782 2142 2785 2148
rect 2774 1892 2777 1978
rect 2762 1848 2766 1851
rect 2782 1802 2785 2078
rect 2790 1922 2793 2148
rect 2798 1972 2801 2328
rect 2822 2222 2825 2478
rect 2838 2352 2841 2558
rect 2846 2492 2849 2668
rect 2854 2462 2857 2698
rect 2862 2652 2865 2668
rect 2862 2532 2865 2558
rect 2870 2512 2873 2558
rect 2878 2522 2881 2908
rect 2904 2903 2906 2907
rect 2910 2903 2913 2907
rect 2918 2903 2920 2907
rect 2886 2572 2889 2888
rect 2926 2882 2929 2918
rect 2914 2788 2918 2791
rect 2926 2732 2929 2878
rect 2904 2703 2906 2707
rect 2910 2703 2913 2707
rect 2918 2703 2920 2707
rect 2898 2668 2902 2671
rect 2894 2582 2897 2648
rect 2902 2642 2905 2668
rect 2926 2622 2929 2728
rect 2894 2542 2897 2578
rect 2866 2478 2870 2481
rect 2878 2462 2881 2508
rect 2904 2503 2906 2507
rect 2910 2503 2913 2507
rect 2918 2503 2920 2507
rect 2854 2342 2857 2348
rect 2830 2332 2833 2338
rect 2818 2148 2825 2151
rect 2822 2142 2825 2148
rect 2822 2102 2825 2118
rect 2806 2092 2809 2098
rect 2814 1832 2817 2078
rect 2758 1762 2761 1768
rect 2754 1748 2758 1751
rect 2774 1662 2777 1668
rect 2802 1558 2806 1561
rect 2814 1512 2817 1738
rect 2822 1662 2825 2098
rect 2830 2092 2833 2328
rect 2846 2302 2849 2338
rect 2862 2322 2865 2338
rect 2870 2332 2873 2338
rect 2846 2282 2849 2298
rect 2846 2152 2849 2258
rect 2878 2222 2881 2458
rect 2866 2128 2870 2131
rect 2830 2062 2833 2078
rect 2846 1992 2849 2008
rect 2838 1882 2841 1988
rect 2854 1822 2857 2028
rect 2870 1912 2873 1968
rect 2878 1932 2881 2128
rect 2894 2112 2897 2348
rect 2926 2312 2929 2318
rect 2904 2303 2906 2307
rect 2910 2303 2913 2307
rect 2918 2303 2920 2307
rect 2894 2042 2897 2108
rect 2904 2103 2906 2107
rect 2910 2103 2913 2107
rect 2918 2103 2920 2107
rect 2926 2102 2929 2138
rect 2890 1918 2894 1921
rect 2904 1903 2906 1907
rect 2910 1903 2913 1907
rect 2918 1903 2920 1907
rect 2926 1902 2929 2068
rect 2934 2022 2937 2688
rect 2942 2152 2945 3518
rect 2958 3452 2961 3458
rect 2966 3252 2969 3268
rect 2974 2962 2977 3588
rect 3334 3552 3337 3588
rect 3150 3532 3153 3548
rect 3210 3538 3214 3541
rect 3322 3538 3326 3541
rect 3014 3452 3017 3458
rect 3006 3282 3009 3318
rect 3014 3271 3017 3378
rect 3010 3268 3017 3271
rect 3014 3072 3017 3258
rect 3022 2762 3025 3358
rect 3038 3292 3041 3528
rect 3030 3022 3033 3128
rect 3062 3062 3065 3268
rect 3150 3252 3153 3528
rect 3262 3511 3265 3528
rect 3258 3508 3265 3511
rect 3202 3448 3206 3451
rect 3174 3332 3177 3338
rect 3174 3272 3177 3278
rect 3138 3158 3142 3161
rect 3118 3112 3121 3128
rect 3046 2682 3049 2848
rect 2998 2552 3001 2578
rect 2942 2132 2945 2148
rect 2950 2122 2953 2458
rect 2986 2448 2990 2451
rect 3022 2442 3025 2498
rect 3054 2442 3057 2978
rect 3118 2972 3121 3048
rect 3062 2472 3065 2638
rect 3070 2482 3073 2528
rect 3070 2472 3073 2478
rect 2990 2392 2993 2398
rect 2958 2142 2961 2358
rect 2990 2261 2993 2388
rect 2998 2342 3001 2348
rect 2986 2258 2993 2261
rect 2962 2128 2966 2131
rect 2934 1912 2937 1968
rect 2962 1928 2966 1931
rect 2974 1922 2977 1938
rect 2918 1872 2921 1878
rect 2870 1762 2873 1858
rect 2862 1752 2865 1758
rect 2870 1742 2873 1748
rect 2846 1682 2849 1688
rect 2842 1668 2846 1671
rect 2830 1542 2833 1598
rect 2854 1501 2857 1508
rect 2870 1502 2873 1518
rect 2854 1498 2862 1501
rect 2758 1452 2761 1478
rect 2694 1412 2697 1438
rect 2798 1412 2801 1428
rect 2794 1358 2801 1361
rect 2630 732 2633 848
rect 2654 802 2657 848
rect 2662 662 2665 938
rect 2678 862 2681 868
rect 2686 832 2689 938
rect 2694 862 2697 1088
rect 2706 1048 2710 1051
rect 2702 782 2705 948
rect 2710 872 2713 908
rect 2698 748 2702 751
rect 2678 732 2681 748
rect 2686 732 2689 748
rect 2590 482 2593 548
rect 2622 542 2625 608
rect 2690 558 2694 561
rect 2510 232 2513 248
rect 2518 242 2521 248
rect 2510 12 2513 228
rect 2558 132 2561 468
rect 2626 438 2630 441
rect 2566 352 2569 368
rect 2574 312 2577 428
rect 2630 392 2633 438
rect 2646 352 2649 428
rect 2598 322 2601 338
rect 2654 332 2657 468
rect 2686 438 2694 441
rect 2590 272 2593 298
rect 2594 268 2598 271
rect 2606 72 2609 268
rect 2686 162 2689 438
rect 2702 352 2705 638
rect 2718 602 2721 958
rect 2726 592 2729 1128
rect 2742 962 2745 1188
rect 2750 1092 2753 1128
rect 2758 1072 2761 1258
rect 2782 1172 2785 1268
rect 2754 1048 2758 1051
rect 2790 1042 2793 1338
rect 2798 1332 2801 1358
rect 2806 1172 2809 1448
rect 2826 1288 2830 1291
rect 2806 1072 2809 1128
rect 2806 1062 2809 1068
rect 2742 952 2745 958
rect 2762 948 2766 951
rect 2742 582 2745 938
rect 2766 892 2769 898
rect 2750 872 2753 878
rect 2766 772 2769 888
rect 2782 858 2790 861
rect 2710 322 2713 548
rect 2718 462 2721 538
rect 2742 462 2745 538
rect 2734 352 2737 458
rect 2722 348 2726 351
rect 2706 168 2710 171
rect 2722 148 2726 151
rect 2690 138 2694 141
rect 2742 72 2745 378
rect 2750 362 2753 768
rect 2774 692 2777 858
rect 2782 672 2785 858
rect 2798 822 2801 988
rect 2806 952 2809 988
rect 2814 872 2817 1068
rect 2830 962 2833 1048
rect 2838 1032 2841 1478
rect 2850 1468 2854 1471
rect 2886 1382 2889 1708
rect 2904 1703 2906 1707
rect 2910 1703 2913 1707
rect 2918 1703 2920 1707
rect 2904 1503 2906 1507
rect 2910 1503 2913 1507
rect 2918 1503 2920 1507
rect 2846 1372 2849 1378
rect 2870 1358 2878 1361
rect 2862 1072 2865 1338
rect 2870 1332 2873 1358
rect 2930 1308 2937 1311
rect 2904 1303 2906 1307
rect 2910 1303 2913 1307
rect 2918 1303 2920 1307
rect 2934 1292 2937 1308
rect 2942 1182 2945 1858
rect 2950 1452 2953 1768
rect 2966 1722 2969 1908
rect 2982 1752 2985 1858
rect 2958 1702 2961 1718
rect 2950 1262 2953 1448
rect 2958 1372 2961 1388
rect 2962 1328 2966 1331
rect 2838 961 2841 1028
rect 2838 958 2846 961
rect 2830 882 2833 948
rect 2838 832 2841 948
rect 2854 882 2857 1068
rect 2866 1038 2870 1041
rect 2866 948 2870 951
rect 2846 872 2849 878
rect 2854 852 2857 868
rect 2822 702 2825 828
rect 2838 792 2841 828
rect 2774 642 2777 648
rect 2782 638 2790 641
rect 2766 582 2769 608
rect 2774 602 2777 608
rect 2774 522 2777 558
rect 2782 382 2785 638
rect 2798 631 2801 638
rect 2790 628 2801 631
rect 2790 492 2793 628
rect 2806 612 2809 688
rect 2822 572 2825 598
rect 2802 538 2806 541
rect 2790 432 2793 438
rect 2750 342 2753 348
rect 2790 342 2793 398
rect 2806 302 2809 518
rect 2822 491 2825 518
rect 2818 488 2825 491
rect 2814 458 2822 461
rect 2814 192 2817 458
rect 2830 332 2833 758
rect 2854 732 2857 748
rect 2862 712 2865 928
rect 2870 862 2873 898
rect 2878 882 2881 1148
rect 2904 1103 2906 1107
rect 2910 1103 2913 1107
rect 2918 1103 2920 1107
rect 2934 1102 2937 1138
rect 2942 1112 2945 1168
rect 2950 1162 2953 1198
rect 2958 1122 2961 1328
rect 2966 1192 2969 1258
rect 2982 1252 2985 1748
rect 2990 1732 2993 2038
rect 2998 1872 3001 2188
rect 3006 1952 3009 2018
rect 3022 1952 3025 2368
rect 3030 2192 3033 2348
rect 3062 2342 3065 2468
rect 3078 2402 3081 2648
rect 3038 2262 3041 2268
rect 3054 2262 3057 2288
rect 3038 1942 3041 2238
rect 3086 2182 3089 2768
rect 3114 2678 3118 2681
rect 3102 2562 3105 2618
rect 3126 2542 3129 2978
rect 3118 2492 3121 2538
rect 3114 2418 3118 2421
rect 2990 1692 2993 1708
rect 2998 1692 3001 1868
rect 3006 1672 3009 1678
rect 3022 1492 3025 1808
rect 3010 1468 3014 1471
rect 2990 1292 2993 1298
rect 2986 1228 2990 1231
rect 2966 1152 2969 1188
rect 2998 1132 3001 1458
rect 3006 1272 3009 1408
rect 3014 1382 3017 1408
rect 3006 1232 3009 1268
rect 2854 642 2857 698
rect 2846 562 2849 608
rect 2838 322 2841 478
rect 2854 472 2857 558
rect 2862 502 2865 538
rect 2854 452 2857 458
rect 2854 412 2857 438
rect 2862 372 2865 488
rect 2870 462 2873 678
rect 2878 422 2881 638
rect 2878 412 2881 418
rect 2850 348 2857 351
rect 2854 342 2857 348
rect 2838 142 2841 218
rect 2854 52 2857 338
rect 2862 272 2865 368
rect 2870 282 2873 348
rect 2870 262 2873 278
rect 2886 151 2889 1058
rect 2894 732 2897 908
rect 2904 903 2906 907
rect 2910 903 2913 907
rect 2918 903 2920 907
rect 2906 868 2910 871
rect 2918 862 2921 868
rect 2902 812 2905 838
rect 2902 752 2905 758
rect 2926 752 2929 968
rect 2894 622 2897 728
rect 2904 703 2906 707
rect 2910 703 2913 707
rect 2918 703 2920 707
rect 2906 638 2913 641
rect 2910 562 2913 638
rect 2926 572 2929 708
rect 2934 572 2937 998
rect 2958 971 2961 1028
rect 2954 968 2961 971
rect 2974 952 2977 958
rect 2966 932 2969 948
rect 2946 868 2950 871
rect 2958 771 2961 848
rect 2958 768 2966 771
rect 2946 728 2950 731
rect 2966 702 2969 768
rect 2950 602 2953 698
rect 2934 552 2937 568
rect 2894 512 2897 518
rect 2904 503 2906 507
rect 2910 503 2913 507
rect 2918 503 2920 507
rect 2926 502 2929 528
rect 2930 458 2934 461
rect 2950 461 2953 598
rect 2966 561 2969 668
rect 2962 558 2969 561
rect 2950 458 2958 461
rect 2966 402 2969 558
rect 2974 461 2977 868
rect 2982 842 2985 1038
rect 2990 982 2993 1068
rect 3014 1062 3017 1088
rect 2982 792 2985 808
rect 2990 752 2993 978
rect 2982 732 2985 738
rect 2998 692 3001 948
rect 3006 922 3009 938
rect 3006 872 3009 878
rect 3006 682 3009 838
rect 3014 782 3017 1058
rect 3022 782 3025 1098
rect 3030 1022 3033 1158
rect 3038 1112 3041 1898
rect 3046 1642 3049 2048
rect 3054 1952 3057 2168
rect 3078 2138 3086 2141
rect 3078 2092 3081 2138
rect 3066 1948 3070 1951
rect 3054 1902 3057 1918
rect 3046 1572 3049 1638
rect 3046 1132 3049 1568
rect 3054 1422 3057 1718
rect 3062 1522 3065 1808
rect 3070 1752 3073 1948
rect 3070 1682 3073 1748
rect 3078 1712 3081 2088
rect 3094 2082 3097 2318
rect 3118 2282 3121 2368
rect 3134 2352 3137 2478
rect 3110 2122 3113 2178
rect 3094 1932 3097 2078
rect 3110 2061 3113 2118
rect 3106 2058 3113 2061
rect 3126 2042 3129 2058
rect 3126 1942 3129 2038
rect 3142 1992 3145 3008
rect 3158 2962 3161 3168
rect 3182 3082 3185 3378
rect 3190 2982 3193 3448
rect 3262 3422 3265 3438
rect 3198 3112 3201 3388
rect 3270 3362 3273 3378
rect 3278 3322 3281 3418
rect 3286 3352 3289 3408
rect 3174 2762 3177 2938
rect 3206 2892 3209 3058
rect 3270 2992 3273 3318
rect 3286 3032 3289 3188
rect 3294 2902 3297 3408
rect 3408 3403 3410 3407
rect 3414 3403 3417 3407
rect 3422 3403 3424 3407
rect 3342 3372 3345 3388
rect 3374 3382 3377 3398
rect 3418 3358 3425 3361
rect 3422 3342 3425 3358
rect 3302 2942 3305 3098
rect 3198 2772 3201 2888
rect 3178 2658 3182 2661
rect 3150 2472 3153 2568
rect 3174 2552 3177 2568
rect 3158 2142 3161 2478
rect 3190 2322 3193 2678
rect 3166 2272 3169 2278
rect 3198 2262 3201 2368
rect 3206 2352 3209 2558
rect 3214 2532 3217 2658
rect 3238 2562 3241 2778
rect 3278 2751 3281 2898
rect 3274 2748 3281 2751
rect 3274 2718 3278 2721
rect 3234 2558 3238 2561
rect 3214 2372 3217 2508
rect 3222 2492 3225 2508
rect 3234 2488 3238 2491
rect 3246 2482 3249 2638
rect 3262 2602 3265 2618
rect 3254 2492 3257 2538
rect 3262 2491 3265 2598
rect 3262 2488 3270 2491
rect 3270 2452 3273 2468
rect 3218 2308 3222 2311
rect 3206 2262 3209 2268
rect 3270 2262 3273 2388
rect 3278 2282 3281 2528
rect 3222 2112 3225 2208
rect 3086 1902 3089 1928
rect 3102 1832 3105 1858
rect 3086 1612 3089 1668
rect 3070 1608 3078 1611
rect 3070 1592 3073 1608
rect 3070 1512 3073 1518
rect 3062 1282 3065 1428
rect 3086 1321 3089 1558
rect 3086 1318 3094 1321
rect 3086 1312 3089 1318
rect 3086 1262 3089 1308
rect 3046 1062 3049 1128
rect 3070 1062 3073 1138
rect 3050 1058 3057 1061
rect 3038 1022 3041 1048
rect 3038 981 3041 1008
rect 3034 978 3041 981
rect 3018 768 3025 771
rect 3002 658 3009 661
rect 3006 612 3009 658
rect 2998 572 3001 578
rect 2974 458 2982 461
rect 3022 432 3025 768
rect 2922 348 2926 351
rect 2894 302 2897 328
rect 2990 322 2993 378
rect 3014 352 3017 388
rect 2904 303 2906 307
rect 2910 303 2913 307
rect 2918 303 2920 307
rect 2990 301 2993 318
rect 2986 298 2993 301
rect 3006 262 3009 268
rect 2922 178 2926 181
rect 2974 152 2977 188
rect 3006 161 3009 178
rect 3002 158 3009 161
rect 2886 148 2894 151
rect 3014 142 3017 348
rect 3022 292 3025 398
rect 3030 312 3033 898
rect 3038 662 3041 818
rect 3046 732 3049 1018
rect 3054 772 3057 1058
rect 3062 952 3065 958
rect 3070 941 3073 998
rect 3066 938 3073 941
rect 3070 882 3073 928
rect 3070 832 3073 858
rect 3054 752 3057 768
rect 3038 452 3041 658
rect 3062 342 3065 728
rect 3078 722 3081 1248
rect 3086 972 3089 1118
rect 3094 892 3097 1088
rect 3102 1052 3105 1708
rect 3110 1482 3113 1498
rect 3110 1372 3113 1398
rect 3110 1122 3113 1328
rect 3086 732 3089 878
rect 3110 861 3113 1108
rect 3106 858 3113 861
rect 3118 992 3121 1858
rect 3126 1742 3129 1778
rect 3134 1662 3137 1958
rect 3158 1942 3161 1948
rect 3166 1942 3169 1978
rect 3150 1842 3153 1938
rect 3134 1578 3142 1581
rect 3126 1562 3129 1568
rect 3126 1132 3129 1418
rect 3134 1382 3137 1578
rect 3150 1452 3153 1828
rect 3158 1712 3161 1768
rect 3166 1752 3169 1908
rect 3190 1762 3193 1868
rect 3222 1772 3225 1898
rect 3238 1802 3241 2108
rect 3238 1732 3241 1788
rect 3158 1652 3161 1708
rect 3230 1702 3233 1728
rect 3238 1671 3241 1728
rect 3234 1668 3241 1671
rect 3162 1478 3166 1481
rect 3174 1472 3177 1668
rect 3134 1322 3137 1328
rect 3142 1281 3145 1298
rect 3138 1278 3145 1281
rect 3134 1042 3137 1128
rect 3106 728 3110 731
rect 3094 662 3097 668
rect 3118 662 3121 988
rect 3138 978 3142 981
rect 3150 962 3153 1398
rect 3158 1322 3161 1458
rect 3174 1312 3177 1468
rect 3166 1032 3169 1258
rect 3158 972 3161 1018
rect 3126 772 3129 948
rect 3154 868 3158 871
rect 3074 538 3078 541
rect 3022 252 3025 288
rect 3070 191 3073 498
rect 3102 492 3105 628
rect 3122 598 3126 601
rect 3118 582 3121 588
rect 3110 472 3113 508
rect 3126 282 3129 328
rect 3070 188 3078 191
rect 3034 138 3038 141
rect 2904 103 2906 107
rect 2910 103 2913 107
rect 2918 103 2920 107
rect 3134 102 3137 428
rect 3142 102 3145 818
rect 3166 712 3169 998
rect 3162 658 3166 661
rect 3174 652 3177 1298
rect 3182 1212 3185 1248
rect 3182 932 3185 1208
rect 3190 1132 3193 1588
rect 3206 1352 3209 1418
rect 3190 1092 3193 1128
rect 3198 1122 3201 1158
rect 3206 1152 3209 1348
rect 3214 1282 3217 1488
rect 3222 1332 3225 1568
rect 3230 1532 3233 1538
rect 3238 1532 3241 1638
rect 3246 1562 3249 1928
rect 3254 1908 3262 1911
rect 3254 1842 3257 1908
rect 3270 1882 3273 2218
rect 3278 1902 3281 2278
rect 3286 1942 3289 2708
rect 3310 2142 3313 3068
rect 3318 2962 3321 3258
rect 3374 3252 3377 3258
rect 3408 3203 3410 3207
rect 3414 3203 3417 3207
rect 3422 3203 3424 3207
rect 3346 3158 3350 3161
rect 3398 3038 3406 3041
rect 3330 2948 3334 2951
rect 3342 2851 3345 2978
rect 3378 2948 3382 2951
rect 3390 2852 3393 2958
rect 3342 2848 3350 2851
rect 3398 2712 3401 3038
rect 3408 3003 3410 3007
rect 3414 3003 3417 3007
rect 3422 3003 3424 3007
rect 3470 2951 3473 2978
rect 3466 2948 3473 2951
rect 3486 2892 3489 3538
rect 3510 3072 3513 3468
rect 3534 3442 3537 3568
rect 3610 3548 3614 3551
rect 3650 3538 3654 3541
rect 3598 3522 3601 3528
rect 3518 3362 3521 3368
rect 3542 3262 3545 3408
rect 3550 3252 3553 3278
rect 3506 2968 3510 2971
rect 3414 2822 3417 2828
rect 3408 2803 3410 2807
rect 3414 2803 3417 2807
rect 3422 2803 3424 2807
rect 3334 2262 3337 2568
rect 3346 2448 3350 2451
rect 3302 2072 3305 2078
rect 3294 2062 3297 2068
rect 3294 2022 3297 2048
rect 3302 1952 3305 1958
rect 3270 1861 3273 1878
rect 3266 1858 3273 1861
rect 3270 1822 3273 1848
rect 3270 1552 3273 1798
rect 3278 1732 3281 1898
rect 3286 1762 3289 1938
rect 3310 1902 3313 2128
rect 3318 2112 3321 2258
rect 3326 2122 3329 2128
rect 3322 2068 3326 2071
rect 3326 1972 3329 2068
rect 3342 1901 3345 2298
rect 3350 2112 3353 2428
rect 3358 2332 3361 2378
rect 3374 2092 3377 2708
rect 3408 2603 3410 2607
rect 3414 2603 3417 2607
rect 3422 2603 3424 2607
rect 3398 2591 3401 2598
rect 3398 2588 3409 2591
rect 3406 2532 3409 2588
rect 3414 2572 3417 2578
rect 3382 2402 3385 2528
rect 3394 2478 3398 2481
rect 3394 2468 3398 2471
rect 3438 2442 3441 2858
rect 3408 2403 3410 2407
rect 3414 2403 3417 2407
rect 3422 2403 3424 2407
rect 3446 2362 3449 2788
rect 3494 2602 3497 2958
rect 3494 2542 3497 2598
rect 3482 2468 3486 2471
rect 3434 2278 3438 2281
rect 3408 2203 3410 2207
rect 3414 2203 3417 2207
rect 3422 2203 3424 2207
rect 3398 2142 3401 2198
rect 3370 2078 3374 2081
rect 3354 2058 3358 2061
rect 3374 2052 3377 2058
rect 3342 1898 3353 1901
rect 3230 1252 3233 1528
rect 3238 1492 3241 1518
rect 3262 1482 3265 1528
rect 3190 942 3193 1088
rect 3182 722 3185 808
rect 3198 672 3201 1058
rect 3206 742 3209 858
rect 3186 558 3190 561
rect 3158 532 3161 558
rect 3206 552 3209 658
rect 3214 562 3217 1118
rect 3222 802 3225 1028
rect 3230 972 3233 1198
rect 3238 1172 3241 1238
rect 3174 422 3177 548
rect 3214 452 3217 558
rect 3150 262 3153 368
rect 3214 362 3217 448
rect 3158 172 3161 358
rect 3222 342 3225 478
rect 3174 272 3177 318
rect 3186 278 3190 281
rect 3162 148 3166 151
rect 3138 78 3142 81
rect 3230 72 3233 778
rect 3238 112 3241 1158
rect 3246 1092 3249 1368
rect 3246 742 3249 958
rect 3254 762 3257 948
rect 3270 942 3273 1328
rect 3278 1142 3281 1728
rect 3302 1622 3305 1848
rect 3310 1682 3313 1898
rect 3342 1862 3345 1888
rect 3338 1858 3342 1861
rect 3318 1662 3321 1668
rect 3286 1402 3289 1558
rect 3350 1552 3353 1898
rect 3366 1861 3369 2028
rect 3408 2003 3410 2007
rect 3414 2003 3417 2007
rect 3422 2003 3424 2007
rect 3382 1882 3385 1988
rect 3390 1962 3393 1988
rect 3366 1858 3374 1861
rect 3310 1512 3313 1538
rect 3350 1512 3353 1528
rect 3298 1508 3302 1511
rect 3330 1508 3334 1511
rect 3374 1452 3377 1858
rect 3398 1842 3401 1998
rect 3414 1912 3417 1928
rect 3386 1838 3390 1841
rect 3382 1542 3385 1768
rect 3322 1378 3326 1381
rect 3318 1342 3321 1348
rect 3266 928 3270 931
rect 3262 842 3265 928
rect 3254 642 3257 758
rect 3278 672 3281 1138
rect 3286 1062 3289 1288
rect 3310 1061 3313 1278
rect 3318 1152 3321 1338
rect 3334 1292 3337 1348
rect 3342 1272 3345 1358
rect 3374 1342 3377 1358
rect 3358 1292 3361 1318
rect 3358 1192 3361 1258
rect 3390 1152 3393 1818
rect 3408 1803 3410 1807
rect 3414 1803 3417 1807
rect 3422 1803 3424 1807
rect 3430 1752 3433 2188
rect 3442 2058 3446 2061
rect 3438 1962 3441 2018
rect 3438 1932 3441 1958
rect 3446 1942 3449 1978
rect 3434 1728 3438 1731
rect 3398 1682 3401 1688
rect 3326 1092 3329 1148
rect 3306 1058 3313 1061
rect 3294 902 3297 988
rect 3302 882 3305 968
rect 3326 882 3329 998
rect 3294 732 3297 878
rect 3334 742 3337 1138
rect 3386 1128 3390 1131
rect 3354 1068 3361 1071
rect 3358 1062 3361 1068
rect 3294 702 3297 718
rect 3290 688 3294 691
rect 3278 502 3281 528
rect 3270 322 3273 498
rect 3278 332 3281 498
rect 3286 262 3289 508
rect 3302 452 3305 738
rect 3322 718 3326 721
rect 3310 602 3313 608
rect 3318 412 3321 708
rect 3334 652 3337 718
rect 3294 162 3297 218
rect 3294 142 3297 158
rect 3318 62 3321 118
rect 3334 82 3337 358
rect 3342 282 3345 488
rect 3350 272 3353 1048
rect 3358 112 3361 918
rect 3366 782 3369 958
rect 3382 882 3385 888
rect 3378 718 3382 721
rect 3398 691 3401 1658
rect 3408 1603 3410 1607
rect 3414 1603 3417 1607
rect 3422 1603 3424 1607
rect 3446 1582 3449 1918
rect 3454 1472 3457 2438
rect 3462 2392 3465 2418
rect 3478 2372 3481 2448
rect 3494 2332 3497 2518
rect 3462 2282 3465 2288
rect 3462 2052 3465 2078
rect 3462 1472 3465 1748
rect 3408 1403 3410 1407
rect 3414 1403 3417 1407
rect 3422 1403 3424 1407
rect 3422 1272 3425 1368
rect 3408 1203 3410 1207
rect 3414 1203 3417 1207
rect 3422 1203 3424 1207
rect 3426 1118 3433 1121
rect 3430 1092 3433 1118
rect 3426 1068 3430 1071
rect 3408 1003 3410 1007
rect 3414 1003 3417 1007
rect 3422 1003 3424 1007
rect 3406 832 3409 878
rect 3408 803 3410 807
rect 3414 803 3417 807
rect 3422 803 3424 807
rect 3390 688 3401 691
rect 3366 552 3369 678
rect 3366 152 3369 528
rect 3382 522 3385 628
rect 3354 68 3358 71
rect 3366 61 3369 148
rect 3390 62 3393 688
rect 3398 582 3401 678
rect 3408 603 3410 607
rect 3414 603 3417 607
rect 3422 603 3424 607
rect 3430 562 3433 608
rect 3418 528 3425 531
rect 3422 512 3425 528
rect 3430 462 3433 548
rect 3438 532 3441 1468
rect 3462 1462 3465 1468
rect 3454 1432 3457 1458
rect 3446 882 3449 1338
rect 3462 1102 3465 1318
rect 3454 812 3457 1048
rect 3450 758 3454 761
rect 3408 403 3410 407
rect 3414 403 3417 407
rect 3422 403 3424 407
rect 3408 203 3410 207
rect 3414 203 3417 207
rect 3422 203 3424 207
rect 3418 138 3422 141
rect 3430 92 3433 458
rect 3446 212 3449 748
rect 3462 732 3465 1068
rect 3454 682 3457 728
rect 3454 482 3457 588
rect 3462 532 3465 538
rect 3462 361 3465 378
rect 3458 358 3465 361
rect 3470 302 3473 2248
rect 3478 1882 3481 1888
rect 3486 1602 3489 2088
rect 3486 1582 3489 1588
rect 3478 1212 3481 1548
rect 3486 1392 3489 1468
rect 3478 1042 3481 1158
rect 3486 1072 3489 1268
rect 3478 962 3481 968
rect 3486 962 3489 1048
rect 3478 822 3481 848
rect 3486 822 3489 938
rect 3486 442 3489 528
rect 3494 132 3497 2328
rect 3502 1342 3505 2738
rect 3510 2672 3513 2938
rect 3518 2762 3521 2768
rect 3526 2722 3529 3158
rect 3534 3082 3537 3238
rect 3534 3052 3537 3078
rect 3534 2732 3537 3038
rect 3558 3012 3561 3518
rect 3570 3478 3574 3481
rect 3510 2552 3513 2578
rect 3510 1932 3513 1958
rect 3518 1761 3521 2718
rect 3526 2082 3529 2698
rect 3542 2692 3545 2878
rect 3550 2652 3553 2928
rect 3570 2868 3577 2871
rect 3558 2702 3561 2768
rect 3574 2752 3577 2868
rect 3558 2652 3561 2698
rect 3566 2482 3569 2558
rect 3534 2122 3537 2128
rect 3542 2062 3545 2278
rect 3550 2242 3553 2338
rect 3558 2252 3561 2368
rect 3566 2282 3569 2308
rect 3562 2248 3566 2251
rect 3566 2052 3569 2138
rect 3526 1852 3529 2028
rect 3542 1802 3545 2038
rect 3510 1758 3521 1761
rect 3538 1758 3542 1761
rect 3510 1572 3513 1758
rect 3518 1672 3521 1748
rect 3526 1682 3529 1718
rect 3538 1708 3542 1711
rect 3510 1552 3513 1558
rect 3510 1352 3513 1358
rect 3506 1318 3510 1321
rect 3510 1272 3513 1318
rect 3510 1082 3513 1118
rect 3502 682 3505 1078
rect 3510 1032 3513 1048
rect 3510 952 3513 1028
rect 3510 862 3513 928
rect 3510 622 3513 828
rect 3506 548 3510 551
rect 3506 538 3510 541
rect 3510 502 3513 508
rect 3518 442 3521 1668
rect 3550 1532 3553 2018
rect 3562 1928 3566 1931
rect 3566 1852 3569 1888
rect 3558 1842 3561 1848
rect 3574 1652 3577 2728
rect 3558 1521 3561 1618
rect 3550 1518 3561 1521
rect 3534 1462 3537 1468
rect 3542 1362 3545 1478
rect 3526 1082 3529 1348
rect 3542 1172 3545 1348
rect 3534 1142 3537 1148
rect 3526 1062 3529 1078
rect 3550 1072 3553 1518
rect 3574 1482 3577 1638
rect 3574 1342 3577 1478
rect 3582 1402 3585 3478
rect 3590 3362 3593 3438
rect 3590 3052 3593 3188
rect 3598 3052 3601 3488
rect 3590 2582 3593 2758
rect 3590 2482 3593 2488
rect 3598 2382 3601 2608
rect 3606 2172 3609 3488
rect 3614 3092 3617 3438
rect 3622 3162 3625 3318
rect 3614 2742 3617 3078
rect 3622 3062 3625 3078
rect 3622 2872 3625 2948
rect 3614 2152 3617 2548
rect 3622 2462 3625 2688
rect 3602 2148 3606 2151
rect 3590 1852 3593 1958
rect 3590 1662 3593 1798
rect 3562 1258 3566 1261
rect 3574 1252 3577 1338
rect 3582 1252 3585 1368
rect 3582 1172 3585 1248
rect 3526 952 3529 1058
rect 3546 958 3550 961
rect 3518 332 3521 418
rect 3526 62 3529 948
rect 3546 758 3550 761
rect 3534 412 3537 678
rect 3542 492 3545 748
rect 3558 702 3561 1058
rect 3566 942 3569 968
rect 3558 632 3561 648
rect 3554 548 3558 551
rect 3558 532 3561 538
rect 3554 478 3558 481
rect 3554 348 3558 351
rect 3566 202 3569 938
rect 3574 462 3577 738
rect 3582 712 3585 1158
rect 3590 1122 3593 1648
rect 3598 1492 3601 1788
rect 3598 1352 3601 1458
rect 3606 1442 3609 2138
rect 3614 1942 3617 2148
rect 3622 2142 3625 2418
rect 3622 2032 3625 2058
rect 3614 1392 3617 1488
rect 3622 1452 3625 1838
rect 3598 1252 3601 1348
rect 3614 1332 3617 1358
rect 3590 872 3593 1108
rect 3590 782 3593 868
rect 3590 662 3593 768
rect 3598 752 3601 1248
rect 3606 1082 3609 1288
rect 3622 1262 3625 1438
rect 3630 1412 3633 3468
rect 3630 1262 3633 1368
rect 3606 1032 3609 1068
rect 3606 802 3609 998
rect 3574 272 3577 448
rect 3582 182 3585 588
rect 3598 562 3601 708
rect 3594 328 3598 331
rect 3554 168 3558 171
rect 3574 162 3577 168
rect 3558 152 3561 158
rect 3606 152 3609 798
rect 3614 752 3617 1058
rect 3622 992 3625 1238
rect 3630 1122 3633 1258
rect 3630 962 3633 1118
rect 3638 1002 3641 3448
rect 3650 3438 3654 3441
rect 3646 3102 3649 3348
rect 3654 2882 3657 2958
rect 3650 2748 3654 2751
rect 3646 2522 3649 2718
rect 3654 2642 3657 2648
rect 3646 2122 3649 2518
rect 3654 2061 3657 2488
rect 3662 2242 3665 3548
rect 3722 3528 3726 3531
rect 3670 3432 3673 3438
rect 3670 2951 3673 3418
rect 3678 3342 3681 3388
rect 3670 2948 3678 2951
rect 3670 2422 3673 2918
rect 3686 2512 3689 3458
rect 3694 3362 3697 3368
rect 3694 3262 3697 3358
rect 3694 2942 3697 3088
rect 3702 3082 3705 3458
rect 3710 3102 3713 3528
rect 3718 3342 3721 3478
rect 3718 3232 3721 3338
rect 3726 3092 3729 3378
rect 3706 3078 3710 3081
rect 3670 2062 3673 2408
rect 3678 2102 3681 2488
rect 3694 2372 3697 2938
rect 3686 2282 3689 2288
rect 3694 2262 3697 2358
rect 3702 2292 3705 2878
rect 3694 2162 3697 2258
rect 3654 2058 3665 2061
rect 3654 2042 3657 2048
rect 3646 1762 3649 2038
rect 3646 1722 3649 1758
rect 3646 1612 3649 1708
rect 3646 1432 3649 1598
rect 3654 1552 3657 1888
rect 3646 1372 3649 1428
rect 3654 1362 3657 1548
rect 3650 1348 3654 1351
rect 3646 1162 3649 1328
rect 3622 832 3625 868
rect 3630 851 3633 888
rect 3630 848 3638 851
rect 3614 722 3617 728
rect 3614 272 3617 708
rect 3622 702 3625 728
rect 3622 362 3625 688
rect 3630 592 3633 848
rect 3646 841 3649 1098
rect 3654 892 3657 1278
rect 3662 922 3665 2058
rect 3670 1962 3673 2048
rect 3670 1642 3673 1748
rect 3670 1371 3673 1508
rect 3678 1502 3681 2098
rect 3686 1961 3689 2158
rect 3686 1958 3697 1961
rect 3686 1542 3689 1948
rect 3694 1842 3697 1958
rect 3702 1742 3705 2278
rect 3710 2142 3713 2148
rect 3698 1728 3702 1731
rect 3694 1531 3697 1658
rect 3710 1572 3713 1948
rect 3686 1528 3697 1531
rect 3686 1442 3689 1528
rect 3694 1482 3697 1488
rect 3698 1468 3702 1471
rect 3670 1368 3681 1371
rect 3670 1342 3673 1358
rect 3670 1242 3673 1328
rect 3646 838 3657 841
rect 3638 372 3641 508
rect 3634 358 3638 361
rect 3622 252 3625 328
rect 3630 91 3633 338
rect 3630 88 3638 91
rect 3586 68 3590 71
rect 3366 58 3374 61
rect 3482 58 3486 61
rect 3330 38 3334 41
rect 3386 38 3390 41
rect 3646 32 3649 828
rect 3654 512 3657 838
rect 3662 822 3665 908
rect 3654 492 3657 498
rect 3654 452 3657 478
rect 3662 352 3665 788
rect 3670 722 3673 918
rect 3678 741 3681 1368
rect 3686 1322 3689 1418
rect 3686 1272 3689 1288
rect 3686 1252 3689 1258
rect 3686 832 3689 1238
rect 3694 862 3697 1448
rect 3678 738 3689 741
rect 3670 652 3673 658
rect 3678 642 3681 708
rect 3670 602 3673 638
rect 3670 452 3673 578
rect 3670 362 3673 368
rect 3686 152 3689 738
rect 3678 142 3681 148
rect 3694 72 3697 858
rect 3702 462 3705 1438
rect 3710 1072 3713 1548
rect 3718 1361 3721 2718
rect 3726 2262 3729 2858
rect 3734 2722 3737 3538
rect 3742 3472 3745 3478
rect 3742 2812 3745 3448
rect 3750 3052 3753 3088
rect 3758 2932 3761 3318
rect 3734 2542 3737 2548
rect 3742 2482 3745 2768
rect 3750 2472 3753 2888
rect 3726 1552 3729 2258
rect 3734 2052 3737 2268
rect 3734 2032 3737 2038
rect 3734 1692 3737 1838
rect 3734 1602 3737 1658
rect 3726 1422 3729 1538
rect 3726 1372 3729 1388
rect 3718 1358 3729 1361
rect 3710 732 3713 1018
rect 3710 532 3713 658
rect 3710 392 3713 528
rect 3718 502 3721 1318
rect 3710 342 3713 348
rect 3714 168 3718 171
rect 3718 152 3721 158
rect 3706 128 3710 131
rect 3714 78 3718 81
rect 3726 52 3729 1358
rect 3734 782 3737 1588
rect 3734 222 3737 768
rect 3742 112 3745 2368
rect 3750 1852 3753 2088
rect 3758 1952 3761 2928
rect 3758 1932 3761 1938
rect 3758 1862 3761 1868
rect 3750 1742 3753 1748
rect 3750 1652 3753 1668
rect 3750 1262 3753 1638
rect 3758 1572 3761 1828
rect 3750 1242 3753 1248
rect 3758 1212 3761 1458
rect 3758 772 3761 1188
rect 3758 652 3761 698
rect 3754 338 3758 341
rect 3758 72 3761 78
rect 3766 62 3769 3268
rect 3774 2652 3777 3448
rect 3774 1462 3777 2098
rect 3774 1432 3777 1448
rect 3774 762 3777 1358
rect 3822 332 3825 2548
rect 726 8 734 11
rect 344 3 346 7
rect 350 3 353 7
rect 358 3 360 7
rect 1360 3 1362 7
rect 1366 3 1369 7
rect 1374 3 1376 7
rect 2384 3 2386 7
rect 2390 3 2393 7
rect 2398 3 2400 7
rect 3408 3 3410 7
rect 3414 3 3417 7
rect 3422 3 3424 7
<< m5contact >>
rect 346 3603 350 3607
rect 353 3603 354 3607
rect 354 3603 357 3607
rect 1362 3603 1366 3607
rect 1369 3603 1370 3607
rect 1370 3603 1373 3607
rect 2386 3603 2390 3607
rect 2393 3603 2394 3607
rect 2394 3603 2397 3607
rect 3410 3603 3414 3607
rect 3417 3603 3418 3607
rect 3418 3603 3421 3607
rect 142 3268 146 3272
rect 38 2848 42 2852
rect 118 2848 122 2852
rect 6 1958 10 1962
rect 14 1848 18 1852
rect 6 1658 10 1662
rect 14 1338 18 1342
rect 46 1948 50 1952
rect 134 2748 138 2752
rect 134 2488 138 2492
rect 134 2128 138 2132
rect 190 2438 194 2442
rect 134 1728 138 1732
rect 118 1668 122 1672
rect 94 1628 98 1632
rect 14 1168 18 1172
rect 14 1148 18 1152
rect 22 1068 26 1072
rect 54 1058 58 1062
rect 86 888 90 892
rect 62 728 66 732
rect 86 688 90 692
rect 198 1938 202 1942
rect 174 1318 178 1322
rect 102 728 106 732
rect 174 688 178 692
rect 346 3403 350 3407
rect 353 3403 354 3407
rect 354 3403 357 3407
rect 346 3203 350 3207
rect 353 3203 354 3207
rect 354 3203 357 3207
rect 346 3003 350 3007
rect 353 3003 354 3007
rect 354 3003 357 3007
rect 254 2848 258 2852
rect 346 2803 350 2807
rect 353 2803 354 2807
rect 354 2803 357 2807
rect 346 2603 350 2607
rect 353 2603 354 2607
rect 354 2603 357 2607
rect 374 2638 378 2642
rect 346 2403 350 2407
rect 353 2403 354 2407
rect 354 2403 357 2407
rect 346 2203 350 2207
rect 353 2203 354 2207
rect 354 2203 357 2207
rect 346 2003 350 2007
rect 353 2003 354 2007
rect 354 2003 357 2007
rect 346 1803 350 1807
rect 353 1803 354 1807
rect 354 1803 357 1807
rect 346 1603 350 1607
rect 353 1603 354 1607
rect 354 1603 357 1607
rect 346 1403 350 1407
rect 353 1403 354 1407
rect 354 1403 357 1407
rect 510 3238 514 3242
rect 502 2668 506 2672
rect 478 2628 482 2632
rect 346 1203 350 1207
rect 353 1203 354 1207
rect 354 1203 357 1207
rect 326 1058 330 1062
rect 346 1003 350 1007
rect 353 1003 354 1007
rect 354 1003 357 1007
rect 318 898 322 902
rect 346 803 350 807
rect 353 803 354 807
rect 354 803 357 807
rect 346 603 350 607
rect 353 603 354 607
rect 354 603 357 607
rect 478 1938 482 1942
rect 478 1738 482 1742
rect 542 2468 546 2472
rect 598 3028 602 3032
rect 646 2568 650 2572
rect 670 2988 674 2992
rect 670 2648 674 2652
rect 662 2558 666 2562
rect 646 2368 650 2372
rect 678 2368 682 2372
rect 478 1328 482 1332
rect 526 1658 530 1662
rect 534 1358 538 1362
rect 494 688 498 692
rect 382 488 386 492
rect 346 403 350 407
rect 353 403 354 407
rect 354 403 357 407
rect 534 1138 538 1142
rect 558 1338 562 1342
rect 606 1848 610 1852
rect 558 1168 562 1172
rect 542 898 546 902
rect 542 338 546 342
rect 478 278 482 282
rect 566 878 570 882
rect 654 1738 658 1742
rect 294 268 298 272
rect 346 203 350 207
rect 353 203 354 207
rect 354 203 357 207
rect 510 68 514 72
rect 850 3503 854 3507
rect 857 3503 858 3507
rect 858 3503 861 3507
rect 910 3538 914 3542
rect 774 3418 778 3422
rect 750 2938 754 2942
rect 726 2658 730 2662
rect 726 2638 730 2642
rect 734 2468 738 2472
rect 766 2868 770 2872
rect 766 2858 770 2862
rect 758 2768 762 2772
rect 766 2678 770 2682
rect 850 3303 854 3307
rect 857 3303 858 3307
rect 858 3303 861 3307
rect 850 3103 854 3107
rect 857 3103 858 3107
rect 858 3103 861 3107
rect 790 2868 794 2872
rect 710 1938 714 1942
rect 662 1468 666 1472
rect 662 1388 666 1392
rect 758 2248 762 2252
rect 750 2138 754 2142
rect 734 1948 738 1952
rect 758 1938 762 1942
rect 814 2788 818 2792
rect 830 2778 834 2782
rect 806 2768 810 2772
rect 822 2728 826 2732
rect 798 2688 802 2692
rect 798 2628 802 2632
rect 798 2548 802 2552
rect 894 3038 898 3042
rect 850 2903 854 2907
rect 857 2903 858 2907
rect 858 2903 861 2907
rect 854 2868 858 2872
rect 838 2718 842 2722
rect 850 2703 854 2707
rect 857 2703 858 2707
rect 858 2703 861 2707
rect 982 3478 986 3482
rect 982 3268 986 3272
rect 974 3158 978 3162
rect 950 2988 954 2992
rect 878 2738 882 2742
rect 854 2628 858 2632
rect 850 2503 854 2507
rect 857 2503 858 2507
rect 858 2503 861 2507
rect 838 2468 842 2472
rect 878 2668 882 2672
rect 878 2638 882 2642
rect 894 2778 898 2782
rect 894 2718 898 2722
rect 878 2528 882 2532
rect 910 2548 914 2552
rect 782 1888 786 1892
rect 850 2303 854 2307
rect 857 2303 858 2307
rect 858 2303 861 2307
rect 814 1738 818 1742
rect 774 1718 778 1722
rect 850 2103 854 2107
rect 857 2103 858 2107
rect 858 2103 861 2107
rect 838 1948 842 1952
rect 850 1903 854 1907
rect 857 1903 858 1907
rect 858 1903 861 1907
rect 850 1703 854 1707
rect 857 1703 858 1707
rect 858 1703 861 1707
rect 942 2698 946 2702
rect 998 3168 1002 3172
rect 990 2788 994 2792
rect 974 2688 978 2692
rect 1014 2768 1018 2772
rect 1014 2758 1018 2762
rect 1006 2628 1010 2632
rect 982 2488 986 2492
rect 990 2458 994 2462
rect 998 2348 1002 2352
rect 1038 3048 1042 3052
rect 1030 2658 1034 2662
rect 1118 3338 1122 3342
rect 1022 2558 1026 2562
rect 1118 2848 1122 2852
rect 1126 2788 1130 2792
rect 1166 3468 1170 3472
rect 1150 2758 1154 2762
rect 1086 2688 1090 2692
rect 1094 2538 1098 2542
rect 966 2138 970 2142
rect 830 1518 834 1522
rect 850 1503 854 1507
rect 857 1503 858 1507
rect 858 1503 861 1507
rect 782 1388 786 1392
rect 702 1138 706 1142
rect 654 678 658 682
rect 814 1328 818 1332
rect 790 488 794 492
rect 806 488 810 492
rect 850 1303 854 1307
rect 857 1303 858 1307
rect 858 1303 861 1307
rect 1094 2268 1098 2272
rect 1078 2248 1082 2252
rect 990 1958 994 1962
rect 998 1948 1002 1952
rect 918 1848 922 1852
rect 910 1688 914 1692
rect 926 1718 930 1722
rect 942 1718 946 1722
rect 1134 2448 1138 2452
rect 1126 2168 1130 2172
rect 1294 3518 1298 3522
rect 1182 3278 1186 3282
rect 1230 3048 1234 3052
rect 1254 2968 1258 2972
rect 1222 2958 1226 2962
rect 1246 2938 1250 2942
rect 1182 2818 1186 2822
rect 1158 2158 1162 2162
rect 1198 2448 1202 2452
rect 1214 2468 1218 2472
rect 1214 2438 1218 2442
rect 1174 2088 1178 2092
rect 1150 2058 1154 2062
rect 998 1668 1002 1672
rect 942 1648 946 1652
rect 982 1638 986 1642
rect 850 1103 854 1107
rect 857 1103 858 1107
rect 858 1103 861 1107
rect 894 1068 898 1072
rect 850 903 854 907
rect 857 903 858 907
rect 858 903 861 907
rect 822 718 826 722
rect 850 703 854 707
rect 857 703 858 707
rect 858 703 861 707
rect 850 503 854 507
rect 857 503 858 507
rect 858 503 861 507
rect 910 538 914 542
rect 974 1468 978 1472
rect 966 1308 970 1312
rect 934 1068 938 1072
rect 950 1058 954 1062
rect 1022 1618 1026 1622
rect 1038 1678 1042 1682
rect 1038 1448 1042 1452
rect 998 1148 1002 1152
rect 990 1058 994 1062
rect 1054 1728 1058 1732
rect 1054 1688 1058 1692
rect 1094 1658 1098 1662
rect 1070 1548 1074 1552
rect 1062 1468 1066 1472
rect 1054 1458 1058 1462
rect 1070 1348 1074 1352
rect 1062 1318 1066 1322
rect 1086 1138 1090 1142
rect 1022 1088 1026 1092
rect 1094 1048 1098 1052
rect 1030 868 1034 872
rect 1110 1078 1114 1082
rect 850 303 854 307
rect 857 303 858 307
rect 858 303 861 307
rect 850 103 854 107
rect 857 103 858 107
rect 858 103 861 107
rect 1022 368 1026 372
rect 934 338 938 342
rect 1022 268 1026 272
rect 1070 348 1074 352
rect 1070 178 1074 182
rect 1238 2428 1242 2432
rect 1238 2358 1242 2362
rect 1230 2328 1234 2332
rect 1294 3268 1298 3272
rect 1294 3248 1298 3252
rect 1286 2948 1290 2952
rect 1318 2958 1322 2962
rect 1302 2918 1306 2922
rect 1302 2858 1306 2862
rect 1390 3538 1394 3542
rect 1362 3403 1366 3407
rect 1369 3403 1370 3407
rect 1370 3403 1373 3407
rect 1350 3338 1354 3342
rect 1362 3203 1366 3207
rect 1369 3203 1370 3207
rect 1370 3203 1373 3207
rect 1362 3003 1366 3007
rect 1369 3003 1370 3007
rect 1370 3003 1373 3007
rect 1414 3468 1418 3472
rect 1430 3348 1434 3352
rect 1406 3258 1410 3262
rect 1362 2803 1366 2807
rect 1369 2803 1370 2807
rect 1370 2803 1373 2807
rect 1294 2348 1298 2352
rect 1198 1878 1202 1882
rect 1182 1558 1186 1562
rect 1158 1388 1162 1392
rect 1134 958 1138 962
rect 1150 1248 1154 1252
rect 1310 2228 1314 2232
rect 1362 2603 1366 2607
rect 1369 2603 1370 2607
rect 1370 2603 1373 2607
rect 1362 2403 1366 2407
rect 1369 2403 1370 2407
rect 1370 2403 1373 2407
rect 1358 2258 1362 2262
rect 1362 2203 1366 2207
rect 1369 2203 1370 2207
rect 1370 2203 1373 2207
rect 1362 2003 1366 2007
rect 1369 2003 1370 2007
rect 1370 2003 1373 2007
rect 1278 1948 1282 1952
rect 1206 1638 1210 1642
rect 1166 1218 1170 1222
rect 1158 1038 1162 1042
rect 1158 1028 1162 1032
rect 1102 368 1106 372
rect 1198 1128 1202 1132
rect 1238 1328 1242 1332
rect 1270 1338 1274 1342
rect 1262 1288 1266 1292
rect 1302 1388 1306 1392
rect 1390 2168 1394 2172
rect 1362 1803 1366 1807
rect 1369 1803 1370 1807
rect 1370 1803 1373 1807
rect 1374 1758 1378 1762
rect 1334 1738 1338 1742
rect 1326 1648 1330 1652
rect 1350 1668 1354 1672
rect 1326 1478 1330 1482
rect 1246 1108 1250 1112
rect 1222 1088 1226 1092
rect 1230 1078 1234 1082
rect 1262 1118 1266 1122
rect 1362 1603 1366 1607
rect 1369 1603 1370 1607
rect 1370 1603 1373 1607
rect 1382 1408 1386 1412
rect 1362 1403 1366 1407
rect 1369 1403 1370 1407
rect 1370 1403 1373 1407
rect 1342 1298 1346 1302
rect 1362 1203 1366 1207
rect 1369 1203 1370 1207
rect 1370 1203 1373 1207
rect 1422 3118 1426 3122
rect 1430 2348 1434 2352
rect 1446 2278 1450 2282
rect 1446 2178 1450 2182
rect 1438 2058 1442 2062
rect 1430 1888 1434 1892
rect 1558 3368 1562 3372
rect 1478 2888 1482 2892
rect 1550 3138 1554 3142
rect 1550 2978 1554 2982
rect 1502 2888 1506 2892
rect 1494 2868 1498 2872
rect 1486 2798 1490 2802
rect 1486 2338 1490 2342
rect 1502 2278 1506 2282
rect 1470 1898 1474 1902
rect 1510 2168 1514 2172
rect 1510 1878 1514 1882
rect 1550 2278 1554 2282
rect 1566 2458 1570 2462
rect 1558 2218 1562 2222
rect 1566 1938 1570 1942
rect 1598 3058 1602 3062
rect 1646 3368 1650 3372
rect 1646 3268 1650 3272
rect 1622 3008 1626 3012
rect 1734 3088 1738 3092
rect 1678 3048 1682 3052
rect 1670 2988 1674 2992
rect 1654 2958 1658 2962
rect 1662 2958 1666 2962
rect 1590 2938 1594 2942
rect 1630 2928 1634 2932
rect 1590 2728 1594 2732
rect 1614 2758 1618 2762
rect 1630 2558 1634 2562
rect 1622 2528 1626 2532
rect 1598 2358 1602 2362
rect 1614 2138 1618 2142
rect 1582 1928 1586 1932
rect 1598 1898 1602 1902
rect 1590 1838 1594 1842
rect 1574 1768 1578 1772
rect 1646 2718 1650 2722
rect 1630 1928 1634 1932
rect 1670 2798 1674 2802
rect 1662 2738 1666 2742
rect 1726 2948 1730 2952
rect 1702 2918 1706 2922
rect 1710 2778 1714 2782
rect 1702 2748 1706 2752
rect 1702 2668 1706 2672
rect 1694 2608 1698 2612
rect 1638 1738 1642 1742
rect 1494 1658 1498 1662
rect 1406 1548 1410 1552
rect 1454 1368 1458 1372
rect 1438 1348 1442 1352
rect 1462 1348 1466 1352
rect 1406 1338 1410 1342
rect 1406 1228 1410 1232
rect 1398 1178 1402 1182
rect 1350 1068 1354 1072
rect 1350 1048 1354 1052
rect 1286 1018 1290 1022
rect 1206 918 1210 922
rect 1238 648 1242 652
rect 1230 388 1234 392
rect 1158 288 1162 292
rect 1190 238 1194 242
rect 1142 188 1146 192
rect 1198 158 1202 162
rect 1318 868 1322 872
rect 1362 1003 1366 1007
rect 1369 1003 1370 1007
rect 1370 1003 1373 1007
rect 1438 1148 1442 1152
rect 1438 1088 1442 1092
rect 1470 1118 1474 1122
rect 1462 1068 1466 1072
rect 1414 1048 1418 1052
rect 1422 1008 1426 1012
rect 1550 1458 1554 1462
rect 1526 1128 1530 1132
rect 1502 1058 1506 1062
rect 1486 948 1490 952
rect 1254 458 1258 462
rect 1262 278 1266 282
rect 1286 468 1290 472
rect 1362 803 1366 807
rect 1369 803 1370 807
rect 1370 803 1373 807
rect 1382 788 1386 792
rect 1286 158 1290 162
rect 1362 603 1366 607
rect 1369 603 1370 607
rect 1370 603 1373 607
rect 1366 568 1370 572
rect 1326 548 1330 552
rect 1362 403 1366 407
rect 1369 403 1370 407
rect 1370 403 1373 407
rect 1350 218 1354 222
rect 1362 203 1366 207
rect 1369 203 1370 207
rect 1370 203 1373 207
rect 1406 798 1410 802
rect 1486 838 1490 842
rect 1502 878 1506 882
rect 1510 758 1514 762
rect 1430 518 1434 522
rect 1438 228 1442 232
rect 1398 158 1402 162
rect 1486 578 1490 582
rect 1510 468 1514 472
rect 1486 458 1490 462
rect 1526 1018 1530 1022
rect 1614 1618 1618 1622
rect 1606 1548 1610 1552
rect 1638 1628 1642 1632
rect 1630 1438 1634 1442
rect 1614 1378 1618 1382
rect 1622 1308 1626 1312
rect 1622 1188 1626 1192
rect 1550 998 1554 1002
rect 1614 1108 1618 1112
rect 1574 848 1578 852
rect 1574 768 1578 772
rect 1558 748 1562 752
rect 1542 738 1546 742
rect 1534 598 1538 602
rect 1598 758 1602 762
rect 1606 668 1610 672
rect 1542 548 1546 552
rect 1590 548 1594 552
rect 1518 288 1522 292
rect 1502 278 1506 282
rect 1550 538 1554 542
rect 1646 1138 1650 1142
rect 1638 1068 1642 1072
rect 1670 1868 1674 1872
rect 1686 1938 1690 1942
rect 1678 1798 1682 1802
rect 1662 1258 1666 1262
rect 1678 1418 1682 1422
rect 1702 2178 1706 2182
rect 1734 2768 1738 2772
rect 1742 2768 1746 2772
rect 1734 2748 1738 2752
rect 1742 2728 1746 2732
rect 1782 3288 1786 3292
rect 1806 3538 1810 3542
rect 1798 3168 1802 3172
rect 1726 2538 1730 2542
rect 1718 2378 1722 2382
rect 1718 2318 1722 2322
rect 1734 2288 1738 2292
rect 1734 2188 1738 2192
rect 1734 2068 1738 2072
rect 1766 2818 1770 2822
rect 1758 2548 1762 2552
rect 1798 3018 1802 3022
rect 1790 2808 1794 2812
rect 1882 3503 1886 3507
rect 1889 3503 1890 3507
rect 1890 3503 1893 3507
rect 1870 3478 1874 3482
rect 1846 2938 1850 2942
rect 1838 2918 1842 2922
rect 1790 2648 1794 2652
rect 1782 2488 1786 2492
rect 1766 2208 1770 2212
rect 1782 2268 1786 2272
rect 1814 2738 1818 2742
rect 1814 2728 1818 2732
rect 1882 3303 1886 3307
rect 1889 3303 1890 3307
rect 1890 3303 1893 3307
rect 1894 3258 1898 3262
rect 1918 3348 1922 3352
rect 1882 3103 1886 3107
rect 1889 3103 1890 3107
rect 1890 3103 1893 3107
rect 1902 2918 1906 2922
rect 1882 2903 1886 2907
rect 1889 2903 1890 2907
rect 1890 2903 1893 2907
rect 1862 2828 1866 2832
rect 1830 2698 1834 2702
rect 1822 2678 1826 2682
rect 1814 2548 1818 2552
rect 1830 2548 1834 2552
rect 1774 1938 1778 1942
rect 1798 2038 1802 2042
rect 1790 1818 1794 1822
rect 1718 1428 1722 1432
rect 1702 1368 1706 1372
rect 1702 1178 1706 1182
rect 1734 1178 1738 1182
rect 1726 1168 1730 1172
rect 1670 1108 1674 1112
rect 1662 1068 1666 1072
rect 1662 1058 1666 1062
rect 1638 1038 1642 1042
rect 1646 768 1650 772
rect 1662 998 1666 1002
rect 1726 958 1730 962
rect 1726 828 1730 832
rect 1702 808 1706 812
rect 1854 2538 1858 2542
rect 1870 2758 1874 2762
rect 1882 2703 1886 2707
rect 1889 2703 1890 2707
rect 1890 2703 1893 2707
rect 1870 2688 1874 2692
rect 1886 2608 1890 2612
rect 1882 2503 1886 2507
rect 1889 2503 1890 2507
rect 1890 2503 1893 2507
rect 1838 2368 1842 2372
rect 1854 2338 1858 2342
rect 1846 2268 1850 2272
rect 1882 2303 1886 2307
rect 1889 2303 1890 2307
rect 1890 2303 1893 2307
rect 1854 2248 1858 2252
rect 1926 2638 1930 2642
rect 1910 2498 1914 2502
rect 1910 2488 1914 2492
rect 1998 3538 2002 3542
rect 1974 3518 1978 3522
rect 1958 2968 1962 2972
rect 1942 2708 1946 2712
rect 1846 2178 1850 2182
rect 1902 2178 1906 2182
rect 1830 2028 1834 2032
rect 1838 2018 1842 2022
rect 1854 2148 1858 2152
rect 1926 2148 1930 2152
rect 1882 2103 1886 2107
rect 1889 2103 1890 2107
rect 1890 2103 1893 2107
rect 1958 2678 1962 2682
rect 1934 2058 1938 2062
rect 1806 1918 1810 1922
rect 1926 1978 1930 1982
rect 1882 1903 1886 1907
rect 1889 1903 1890 1907
rect 1890 1903 1893 1907
rect 1870 1728 1874 1732
rect 1882 1703 1886 1707
rect 1889 1703 1890 1707
rect 1890 1703 1893 1707
rect 1926 1718 1930 1722
rect 1910 1678 1914 1682
rect 1882 1503 1886 1507
rect 1889 1503 1890 1507
rect 1890 1503 1893 1507
rect 1974 2968 1978 2972
rect 1998 3048 2002 3052
rect 1982 2778 1986 2782
rect 1990 2768 1994 2772
rect 1966 2388 1970 2392
rect 1990 2258 1994 2262
rect 2014 2978 2018 2982
rect 2006 2928 2010 2932
rect 2038 3078 2042 3082
rect 2062 3048 2066 3052
rect 2054 2978 2058 2982
rect 2030 2748 2034 2752
rect 2030 2318 2034 2322
rect 2006 2298 2010 2302
rect 2014 2228 2018 2232
rect 2022 2208 2026 2212
rect 2022 2188 2026 2192
rect 1958 1848 1962 1852
rect 1958 1558 1962 1562
rect 1942 1488 1946 1492
rect 1878 1478 1882 1482
rect 1910 1448 1914 1452
rect 1942 1438 1946 1442
rect 1886 1408 1890 1412
rect 1870 1358 1874 1362
rect 1886 1358 1890 1362
rect 1838 1318 1842 1322
rect 1838 1298 1842 1302
rect 1766 1018 1770 1022
rect 1774 868 1778 872
rect 1646 588 1650 592
rect 1606 488 1610 492
rect 1550 338 1554 342
rect 1558 298 1562 302
rect 1526 268 1530 272
rect 1534 258 1538 262
rect 1534 248 1538 252
rect 1790 548 1794 552
rect 1582 268 1586 272
rect 1622 218 1626 222
rect 1590 178 1594 182
rect 1654 168 1658 172
rect 1702 268 1706 272
rect 1766 418 1770 422
rect 1774 288 1778 292
rect 1882 1303 1886 1307
rect 1889 1303 1890 1307
rect 1890 1303 1893 1307
rect 1846 1078 1850 1082
rect 1830 1028 1834 1032
rect 1814 988 1818 992
rect 1830 948 1834 952
rect 1882 1103 1886 1107
rect 1889 1103 1890 1107
rect 1890 1103 1893 1107
rect 1870 1008 1874 1012
rect 1870 948 1874 952
rect 1854 938 1858 942
rect 1822 848 1826 852
rect 1814 818 1818 822
rect 1806 678 1810 682
rect 1830 468 1834 472
rect 1882 903 1886 907
rect 1889 903 1890 907
rect 1890 903 1893 907
rect 1894 878 1898 882
rect 1862 798 1866 802
rect 1854 778 1858 782
rect 1870 768 1874 772
rect 1882 703 1886 707
rect 1889 703 1890 707
rect 1890 703 1893 707
rect 1862 688 1866 692
rect 1882 503 1886 507
rect 1889 503 1890 507
rect 1890 503 1893 507
rect 1950 1268 1954 1272
rect 1926 848 1930 852
rect 2030 1878 2034 1882
rect 2006 1788 2010 1792
rect 1966 1188 1970 1192
rect 1958 958 1962 962
rect 1958 918 1962 922
rect 1974 938 1978 942
rect 1918 738 1922 742
rect 1934 738 1938 742
rect 1910 698 1914 702
rect 1926 668 1930 672
rect 1902 488 1906 492
rect 1862 478 1866 482
rect 1990 1718 1994 1722
rect 2214 3418 2218 3422
rect 2078 3058 2082 3062
rect 2054 2878 2058 2882
rect 2070 2868 2074 2872
rect 2126 3318 2130 3322
rect 2126 3088 2130 3092
rect 2118 2978 2122 2982
rect 2134 2978 2138 2982
rect 2126 2938 2130 2942
rect 2134 2908 2138 2912
rect 2070 2858 2074 2862
rect 2166 3048 2170 3052
rect 2390 3538 2394 3542
rect 2270 3528 2274 3532
rect 2238 3518 2242 3522
rect 2270 3458 2274 3462
rect 2294 3318 2298 3322
rect 2222 3158 2226 3162
rect 2198 3128 2202 3132
rect 2230 3108 2234 3112
rect 2238 3048 2242 3052
rect 2214 2968 2218 2972
rect 2206 2918 2210 2922
rect 2158 2858 2162 2862
rect 2062 2558 2066 2562
rect 2046 1688 2050 1692
rect 2110 2658 2114 2662
rect 2126 2618 2130 2622
rect 2070 1798 2074 1802
rect 1998 1308 2002 1312
rect 1990 1028 1994 1032
rect 1958 658 1962 662
rect 1942 468 1946 472
rect 1974 428 1978 432
rect 1870 378 1874 382
rect 1846 338 1850 342
rect 1942 348 1946 352
rect 1882 303 1886 307
rect 1889 303 1890 307
rect 1890 303 1893 307
rect 1910 288 1914 292
rect 1934 278 1938 282
rect 1910 268 1914 272
rect 1950 258 1954 262
rect 1966 258 1970 262
rect 1838 238 1842 242
rect 1882 103 1886 107
rect 1889 103 1890 107
rect 1890 103 1893 107
rect 1662 68 1666 72
rect 2054 1448 2058 1452
rect 2062 1348 2066 1352
rect 2094 2158 2098 2162
rect 2094 2148 2098 2152
rect 2150 2668 2154 2672
rect 2150 2448 2154 2452
rect 2142 2308 2146 2312
rect 2150 2258 2154 2262
rect 2166 2368 2170 2372
rect 2150 2178 2154 2182
rect 2182 2268 2186 2272
rect 2294 3138 2298 3142
rect 2310 3138 2314 3142
rect 2270 3038 2274 3042
rect 2286 3078 2290 3082
rect 2270 2948 2274 2952
rect 2262 2878 2266 2882
rect 2294 3038 2298 3042
rect 2270 2688 2274 2692
rect 2238 2528 2242 2532
rect 2230 2208 2234 2212
rect 2206 2118 2210 2122
rect 2182 2068 2186 2072
rect 2206 2048 2210 2052
rect 2126 1918 2130 1922
rect 2174 1888 2178 1892
rect 2198 1878 2202 1882
rect 2134 1728 2138 1732
rect 2166 1388 2170 1392
rect 2094 1358 2098 1362
rect 2150 1168 2154 1172
rect 2166 1158 2170 1162
rect 2030 1148 2034 1152
rect 2110 1118 2114 1122
rect 2038 1108 2042 1112
rect 2054 1098 2058 1102
rect 2086 1088 2090 1092
rect 2126 1108 2130 1112
rect 2062 938 2066 942
rect 2062 928 2066 932
rect 2062 868 2066 872
rect 2038 838 2042 842
rect 2062 758 2066 762
rect 2022 678 2026 682
rect 2014 458 2018 462
rect 2014 368 2018 372
rect 2062 638 2066 642
rect 2038 568 2042 572
rect 2142 998 2146 1002
rect 2182 1078 2186 1082
rect 2230 2068 2234 2072
rect 2254 2278 2258 2282
rect 2326 3138 2330 3142
rect 2326 3008 2330 3012
rect 2310 2968 2314 2972
rect 2318 2938 2322 2942
rect 2294 2528 2298 2532
rect 2318 2338 2322 2342
rect 2310 2268 2314 2272
rect 2286 2038 2290 2042
rect 2318 1988 2322 1992
rect 2310 1938 2314 1942
rect 2278 1878 2282 1882
rect 2270 1778 2274 1782
rect 2302 1878 2306 1882
rect 2350 2928 2354 2932
rect 2350 2908 2354 2912
rect 2386 3403 2390 3407
rect 2393 3403 2394 3407
rect 2394 3403 2397 3407
rect 2574 3528 2578 3532
rect 2494 3518 2498 3522
rect 2542 3458 2546 3462
rect 2574 3458 2578 3462
rect 2374 3308 2378 3312
rect 2386 3203 2390 3207
rect 2393 3203 2394 3207
rect 2394 3203 2397 3207
rect 2366 3048 2370 3052
rect 2334 2848 2338 2852
rect 2350 2798 2354 2802
rect 2386 3003 2390 3007
rect 2393 3003 2394 3007
rect 2394 3003 2397 3007
rect 2374 2938 2378 2942
rect 2390 2868 2394 2872
rect 2386 2803 2390 2807
rect 2393 2803 2394 2807
rect 2394 2803 2397 2807
rect 2398 2678 2402 2682
rect 2662 3308 2666 3312
rect 2906 3503 2910 3507
rect 2913 3503 2914 3507
rect 2914 3503 2917 3507
rect 2894 3448 2898 3452
rect 2446 3058 2450 3062
rect 2470 3108 2474 3112
rect 2462 3048 2466 3052
rect 2502 2928 2506 2932
rect 2454 2868 2458 2872
rect 2406 2668 2410 2672
rect 2414 2648 2418 2652
rect 2386 2603 2390 2607
rect 2393 2603 2394 2607
rect 2394 2603 2397 2607
rect 2406 2548 2410 2552
rect 2446 2718 2450 2722
rect 2454 2708 2458 2712
rect 2438 2518 2442 2522
rect 2366 2498 2370 2502
rect 2334 2318 2338 2322
rect 2358 2208 2362 2212
rect 2414 2488 2418 2492
rect 2386 2403 2390 2407
rect 2393 2403 2394 2407
rect 2394 2403 2397 2407
rect 2406 2338 2410 2342
rect 2374 2258 2378 2262
rect 2386 2203 2390 2207
rect 2393 2203 2394 2207
rect 2394 2203 2397 2207
rect 2406 2008 2410 2012
rect 2386 2003 2390 2007
rect 2393 2003 2394 2007
rect 2394 2003 2397 2007
rect 2342 1878 2346 1882
rect 2350 1858 2354 1862
rect 2318 1788 2322 1792
rect 2270 1358 2274 1362
rect 2278 1328 2282 1332
rect 2294 1288 2298 1292
rect 2214 1128 2218 1132
rect 2182 1058 2186 1062
rect 2166 1008 2170 1012
rect 2126 978 2130 982
rect 2102 818 2106 822
rect 2126 818 2130 822
rect 2134 788 2138 792
rect 2102 728 2106 732
rect 2102 658 2106 662
rect 2102 648 2106 652
rect 2086 628 2090 632
rect 2206 928 2210 932
rect 2190 898 2194 902
rect 2214 808 2218 812
rect 2214 788 2218 792
rect 2086 568 2090 572
rect 2078 548 2082 552
rect 2046 388 2050 392
rect 2030 348 2034 352
rect 1950 168 1954 172
rect 2158 568 2162 572
rect 2230 648 2234 652
rect 2182 548 2186 552
rect 2134 538 2138 542
rect 2302 1108 2306 1112
rect 2294 1068 2298 1072
rect 2262 848 2266 852
rect 2254 748 2258 752
rect 2254 678 2258 682
rect 2270 678 2274 682
rect 2286 938 2290 942
rect 2286 768 2290 772
rect 2238 618 2242 622
rect 2326 1318 2330 1322
rect 2318 1248 2322 1252
rect 2374 1958 2378 1962
rect 2438 2278 2442 2282
rect 2446 2158 2450 2162
rect 2430 2078 2434 2082
rect 2462 2558 2466 2562
rect 2470 2318 2474 2322
rect 2486 2268 2490 2272
rect 2478 2248 2482 2252
rect 2462 1948 2466 1952
rect 2438 1888 2442 1892
rect 2374 1868 2378 1872
rect 2414 1848 2418 1852
rect 2386 1803 2390 1807
rect 2393 1803 2394 1807
rect 2394 1803 2397 1807
rect 2374 1758 2378 1762
rect 2390 1758 2394 1762
rect 2366 1748 2370 1752
rect 2398 1718 2402 1722
rect 2366 1688 2370 1692
rect 2386 1603 2390 1607
rect 2393 1603 2394 1607
rect 2394 1603 2397 1607
rect 2386 1403 2390 1407
rect 2393 1403 2394 1407
rect 2394 1403 2397 1407
rect 2342 1268 2346 1272
rect 2386 1203 2390 1207
rect 2393 1203 2394 1207
rect 2394 1203 2397 1207
rect 2454 1878 2458 1882
rect 2454 1848 2458 1852
rect 2518 2578 2522 2582
rect 2510 2548 2514 2552
rect 2494 2048 2498 2052
rect 2906 3303 2910 3307
rect 2913 3303 2914 3307
rect 2914 3303 2917 3307
rect 2902 3238 2906 3242
rect 2606 3058 2610 3062
rect 2574 2988 2578 2992
rect 2550 2828 2554 2832
rect 2542 2478 2546 2482
rect 2526 2348 2530 2352
rect 2550 2258 2554 2262
rect 2510 2168 2514 2172
rect 2534 2158 2538 2162
rect 2542 2098 2546 2102
rect 2526 2058 2530 2062
rect 2486 1478 2490 1482
rect 2502 1388 2506 1392
rect 2486 1328 2490 1332
rect 2422 1198 2426 1202
rect 2374 1178 2378 1182
rect 2430 1178 2434 1182
rect 2374 1038 2378 1042
rect 2386 1003 2390 1007
rect 2393 1003 2394 1007
rect 2394 1003 2397 1007
rect 2374 998 2378 1002
rect 2454 1138 2458 1142
rect 2438 1118 2442 1122
rect 2366 928 2370 932
rect 2366 898 2370 902
rect 2386 803 2390 807
rect 2393 803 2394 807
rect 2394 803 2397 807
rect 2350 718 2354 722
rect 2382 718 2386 722
rect 2334 658 2338 662
rect 2310 648 2314 652
rect 2254 558 2258 562
rect 2062 278 2066 282
rect 2334 538 2338 542
rect 2254 458 2258 462
rect 2334 448 2338 452
rect 2174 438 2178 442
rect 2206 388 2210 392
rect 2222 298 2226 302
rect 2230 298 2234 302
rect 2206 278 2210 282
rect 2278 338 2282 342
rect 2190 258 2194 262
rect 2198 178 2202 182
rect 2190 168 2194 172
rect 2446 1048 2450 1052
rect 2510 1318 2514 1322
rect 2582 2888 2586 2892
rect 2590 2538 2594 2542
rect 2598 2378 2602 2382
rect 2662 3028 2666 3032
rect 2662 2858 2666 2862
rect 2646 2598 2650 2602
rect 2638 2368 2642 2372
rect 2622 2338 2626 2342
rect 2606 2308 2610 2312
rect 2622 2268 2626 2272
rect 2686 3118 2690 3122
rect 2702 2938 2706 2942
rect 2906 3103 2910 3107
rect 2913 3103 2914 3107
rect 2914 3103 2917 3107
rect 2694 2868 2698 2872
rect 2686 2648 2690 2652
rect 2686 2638 2690 2642
rect 2822 2958 2826 2962
rect 2790 2878 2794 2882
rect 2710 2378 2714 2382
rect 2766 2708 2770 2712
rect 2774 2648 2778 2652
rect 2758 2638 2762 2642
rect 2590 2088 2594 2092
rect 2606 2088 2610 2092
rect 2582 2078 2586 2082
rect 2590 2058 2594 2062
rect 2534 1858 2538 1862
rect 2590 1488 2594 1492
rect 2606 1488 2610 1492
rect 2590 1478 2594 1482
rect 2566 1368 2570 1372
rect 2478 1168 2482 1172
rect 2494 1158 2498 1162
rect 2486 1138 2490 1142
rect 2470 1108 2474 1112
rect 2518 1118 2522 1122
rect 2478 1098 2482 1102
rect 2470 1068 2474 1072
rect 2494 998 2498 1002
rect 2574 1188 2578 1192
rect 2550 1128 2554 1132
rect 2566 1048 2570 1052
rect 2574 1048 2578 1052
rect 2558 1028 2562 1032
rect 2574 998 2578 1002
rect 2574 968 2578 972
rect 2510 868 2514 872
rect 2478 828 2482 832
rect 2430 798 2434 802
rect 2446 698 2450 702
rect 2414 638 2418 642
rect 2386 603 2390 607
rect 2393 603 2394 607
rect 2394 603 2397 607
rect 2374 598 2378 602
rect 2366 528 2370 532
rect 2366 458 2370 462
rect 2446 548 2450 552
rect 2446 468 2450 472
rect 2382 438 2386 442
rect 2386 403 2390 407
rect 2393 403 2394 407
rect 2394 403 2397 407
rect 2326 338 2330 342
rect 2350 338 2354 342
rect 2374 338 2378 342
rect 2398 258 2402 262
rect 2386 203 2390 207
rect 2393 203 2394 207
rect 2394 203 2397 207
rect 2438 298 2442 302
rect 2494 788 2498 792
rect 2518 768 2522 772
rect 2486 748 2490 752
rect 2502 748 2506 752
rect 2518 728 2522 732
rect 2486 648 2490 652
rect 2462 448 2466 452
rect 2462 408 2466 412
rect 2478 288 2482 292
rect 2454 278 2458 282
rect 2470 268 2474 272
rect 2470 188 2474 192
rect 2526 618 2530 622
rect 2518 598 2522 602
rect 2502 428 2506 432
rect 2510 358 2514 362
rect 2542 488 2546 492
rect 2582 858 2586 862
rect 2670 2038 2674 2042
rect 2686 2038 2690 2042
rect 2654 1858 2658 1862
rect 2630 1818 2634 1822
rect 2646 1658 2650 1662
rect 2598 1068 2602 1072
rect 2598 1058 2602 1062
rect 2678 1808 2682 1812
rect 2670 1738 2674 1742
rect 2678 1308 2682 1312
rect 2646 1218 2650 1222
rect 2662 1178 2666 1182
rect 2638 1158 2642 1162
rect 2630 958 2634 962
rect 2662 988 2666 992
rect 2638 918 2642 922
rect 2598 898 2602 902
rect 2702 1808 2706 1812
rect 2710 1788 2714 1792
rect 2766 2568 2770 2572
rect 2710 1738 2714 1742
rect 2694 1508 2698 1512
rect 2710 1498 2714 1502
rect 2742 1948 2746 1952
rect 2766 2118 2770 2122
rect 2758 1928 2762 1932
rect 2790 2568 2794 2572
rect 2798 2568 2802 2572
rect 2822 2688 2826 2692
rect 2862 2718 2866 2722
rect 2830 2648 2834 2652
rect 2814 2518 2818 2522
rect 2806 2328 2810 2332
rect 2782 2138 2786 2142
rect 2758 1848 2762 1852
rect 2906 2903 2910 2907
rect 2913 2903 2914 2907
rect 2914 2903 2917 2907
rect 2918 2788 2922 2792
rect 2906 2703 2910 2707
rect 2913 2703 2914 2707
rect 2914 2703 2917 2707
rect 2902 2668 2906 2672
rect 2894 2648 2898 2652
rect 2926 2618 2930 2622
rect 2862 2478 2866 2482
rect 2906 2503 2910 2507
rect 2913 2503 2914 2507
rect 2914 2503 2917 2507
rect 2830 2338 2834 2342
rect 2854 2338 2858 2342
rect 2822 2138 2826 2142
rect 2822 2118 2826 2122
rect 2806 2098 2810 2102
rect 2798 1968 2802 1972
rect 2814 1828 2818 1832
rect 2758 1758 2762 1762
rect 2750 1748 2754 1752
rect 2774 1668 2778 1672
rect 2806 1558 2810 1562
rect 2870 2328 2874 2332
rect 2862 2318 2866 2322
rect 2870 2128 2874 2132
rect 2830 2058 2834 2062
rect 2854 2028 2858 2032
rect 2846 2008 2850 2012
rect 2926 2318 2930 2322
rect 2906 2303 2910 2307
rect 2913 2303 2914 2307
rect 2914 2303 2917 2307
rect 2906 2103 2910 2107
rect 2913 2103 2914 2107
rect 2914 2103 2917 2107
rect 2886 1918 2890 1922
rect 2906 1903 2910 1907
rect 2913 1903 2914 1907
rect 2914 1903 2917 1907
rect 2958 3458 2962 3462
rect 2966 3248 2970 3252
rect 3214 3538 3218 3542
rect 3318 3538 3322 3542
rect 3486 3538 3490 3542
rect 3038 3528 3042 3532
rect 3014 3458 3018 3462
rect 3198 3448 3202 3452
rect 3174 3338 3178 3342
rect 3142 3158 3146 3162
rect 3118 3128 3122 3132
rect 3030 3018 3034 3022
rect 3054 2978 3058 2982
rect 3022 2758 3026 2762
rect 2998 2578 3002 2582
rect 2942 2148 2946 2152
rect 2990 2448 2994 2452
rect 3118 2968 3122 2972
rect 3070 2528 3074 2532
rect 3070 2478 3074 2482
rect 2998 2348 3002 2352
rect 2966 2128 2970 2132
rect 2934 1968 2938 1972
rect 2958 1928 2962 1932
rect 2918 1868 2922 1872
rect 2862 1758 2866 1762
rect 2870 1738 2874 1742
rect 2846 1688 2850 1692
rect 2838 1668 2842 1672
rect 2854 1508 2858 1512
rect 2870 1498 2874 1502
rect 2758 1448 2762 1452
rect 2630 848 2634 852
rect 2654 798 2658 802
rect 2678 858 2682 862
rect 2702 1048 2706 1052
rect 2686 828 2690 832
rect 2710 868 2714 872
rect 2678 748 2682 752
rect 2694 748 2698 752
rect 2702 638 2706 642
rect 2622 608 2626 612
rect 2686 558 2690 562
rect 2526 288 2530 292
rect 2518 238 2522 242
rect 2510 228 2514 232
rect 2630 438 2634 442
rect 2566 368 2570 372
rect 2646 348 2650 352
rect 2598 318 2602 322
rect 2590 268 2594 272
rect 2758 1048 2762 1052
rect 2798 1328 2802 1332
rect 2830 1288 2834 1292
rect 2806 1128 2810 1132
rect 2806 1068 2810 1072
rect 2790 1038 2794 1042
rect 2798 988 2802 992
rect 2806 988 2810 992
rect 2742 958 2746 962
rect 2758 948 2762 952
rect 2766 888 2770 892
rect 2750 878 2754 882
rect 2750 768 2754 772
rect 2742 578 2746 582
rect 2718 538 2722 542
rect 2734 458 2738 462
rect 2718 348 2722 352
rect 2702 168 2706 172
rect 2726 148 2730 152
rect 2694 138 2698 142
rect 2854 1468 2858 1472
rect 2906 1703 2910 1707
rect 2913 1703 2914 1707
rect 2914 1703 2917 1707
rect 2906 1503 2910 1507
rect 2913 1503 2914 1507
rect 2914 1503 2917 1507
rect 2846 1368 2850 1372
rect 2906 1303 2910 1307
rect 2913 1303 2914 1307
rect 2914 1303 2917 1307
rect 2934 1288 2938 1292
rect 2982 1748 2986 1752
rect 2958 1388 2962 1392
rect 2958 1328 2962 1332
rect 2950 1198 2954 1202
rect 2830 948 2834 952
rect 2862 1038 2866 1042
rect 2862 948 2866 952
rect 2846 878 2850 882
rect 2854 848 2858 852
rect 2822 828 2826 832
rect 2838 828 2842 832
rect 2774 648 2778 652
rect 2774 598 2778 602
rect 2766 578 2770 582
rect 2774 558 2778 562
rect 2806 608 2810 612
rect 2822 598 2826 602
rect 2798 538 2802 542
rect 2822 518 2826 522
rect 2790 438 2794 442
rect 2782 378 2786 382
rect 2750 348 2754 352
rect 2822 458 2826 462
rect 2854 728 2858 732
rect 2934 1138 2938 1142
rect 2906 1103 2910 1107
rect 2913 1103 2914 1107
rect 2914 1103 2917 1107
rect 3054 2288 3058 2292
rect 3038 2258 3042 2262
rect 3006 1948 3010 1952
rect 3110 2678 3114 2682
rect 3102 2558 3106 2562
rect 3118 2488 3122 2492
rect 3118 2418 3122 2422
rect 3118 2368 3122 2372
rect 2998 1868 3002 1872
rect 2990 1688 2994 1692
rect 3006 1668 3010 1672
rect 3006 1468 3010 1472
rect 2990 1298 2994 1302
rect 2982 1228 2986 1232
rect 2966 1188 2970 1192
rect 3006 1228 3010 1232
rect 2990 1068 2994 1072
rect 2870 858 2874 862
rect 2854 638 2858 642
rect 2846 608 2850 612
rect 2862 538 2866 542
rect 2854 458 2858 462
rect 2854 438 2858 442
rect 2878 418 2882 422
rect 2862 368 2866 372
rect 2838 138 2842 142
rect 2982 1038 2986 1042
rect 2958 1028 2962 1032
rect 2906 903 2910 907
rect 2913 903 2914 907
rect 2914 903 2917 907
rect 2902 868 2906 872
rect 2918 858 2922 862
rect 2902 808 2906 812
rect 2902 748 2906 752
rect 2906 703 2910 707
rect 2913 703 2914 707
rect 2914 703 2917 707
rect 2894 618 2898 622
rect 2974 958 2978 962
rect 2942 868 2946 872
rect 2942 728 2946 732
rect 2950 698 2954 702
rect 2966 698 2970 702
rect 2966 668 2970 672
rect 2950 598 2954 602
rect 2910 558 2914 562
rect 2894 518 2898 522
rect 2906 503 2910 507
rect 2913 503 2914 507
rect 2914 503 2917 507
rect 2926 458 2930 462
rect 3014 1058 3018 1062
rect 2982 808 2986 812
rect 2982 728 2986 732
rect 3006 918 3010 922
rect 3006 878 3010 882
rect 3078 2088 3082 2092
rect 3070 1948 3074 1952
rect 3054 1918 3058 1922
rect 3110 2178 3114 2182
rect 3270 3358 3274 3362
rect 3190 2978 3194 2982
rect 3410 3403 3414 3407
rect 3417 3403 3418 3407
rect 3418 3403 3421 3407
rect 3422 3338 3426 3342
rect 3174 2658 3178 2662
rect 3150 2568 3154 2572
rect 3166 2278 3170 2282
rect 3270 2718 3274 2722
rect 3238 2558 3242 2562
rect 3230 2488 3234 2492
rect 3262 2598 3266 2602
rect 3254 2488 3258 2492
rect 3270 2448 3274 2452
rect 3270 2388 3274 2392
rect 3222 2308 3226 2312
rect 3206 2258 3210 2262
rect 3270 2218 3274 2222
rect 3166 1978 3170 1982
rect 3126 1938 3130 1942
rect 3102 1858 3106 1862
rect 3086 1668 3090 1672
rect 3070 1588 3074 1592
rect 3070 1518 3074 1522
rect 3062 1428 3066 1432
rect 3062 1278 3066 1282
rect 3038 1108 3042 1112
rect 3038 1048 3042 1052
rect 3038 1008 3042 1012
rect 3022 778 3026 782
rect 3006 608 3010 612
rect 2998 578 3002 582
rect 2918 348 2922 352
rect 2990 318 2994 322
rect 2906 303 2910 307
rect 2913 303 2914 307
rect 2914 303 2917 307
rect 3006 268 3010 272
rect 2918 178 2922 182
rect 3006 178 3010 182
rect 2974 148 2978 152
rect 3062 958 3066 962
rect 3070 928 3074 932
rect 3070 858 3074 862
rect 3086 1118 3090 1122
rect 3110 1478 3114 1482
rect 3110 1118 3114 1122
rect 3126 1778 3130 1782
rect 3158 1938 3162 1942
rect 3150 1838 3154 1842
rect 3126 1568 3130 1572
rect 3158 1768 3162 1772
rect 3238 1798 3242 1802
rect 3230 1728 3234 1732
rect 3238 1728 3242 1732
rect 3158 1708 3162 1712
rect 3166 1478 3170 1482
rect 3190 1588 3194 1592
rect 3134 1328 3138 1332
rect 3142 1298 3146 1302
rect 3134 1038 3138 1042
rect 3118 988 3122 992
rect 3086 728 3090 732
rect 3102 728 3106 732
rect 3134 978 3138 982
rect 3174 1308 3178 1312
rect 3158 1018 3162 1022
rect 3150 868 3154 872
rect 3126 768 3130 772
rect 3094 658 3098 662
rect 3070 538 3074 542
rect 3070 498 3074 502
rect 3022 288 3026 292
rect 3126 598 3130 602
rect 3118 588 3122 592
rect 3110 508 3114 512
rect 3110 468 3114 472
rect 3126 328 3130 332
rect 3038 138 3042 142
rect 2906 103 2910 107
rect 2913 103 2914 107
rect 2914 103 2917 107
rect 3166 708 3170 712
rect 3158 658 3162 662
rect 3182 1248 3186 1252
rect 3206 1418 3210 1422
rect 3374 3248 3378 3252
rect 3410 3203 3414 3207
rect 3417 3203 3418 3207
rect 3418 3203 3421 3207
rect 3342 3158 3346 3162
rect 3326 2948 3330 2952
rect 3374 2948 3378 2952
rect 3410 3003 3414 3007
rect 3417 3003 3418 3007
rect 3418 3003 3421 3007
rect 3470 2978 3474 2982
rect 3606 3548 3610 3552
rect 3646 3538 3650 3542
rect 3598 3518 3602 3522
rect 3518 3368 3522 3372
rect 3502 2968 3506 2972
rect 3414 2818 3418 2822
rect 3410 2803 3414 2807
rect 3417 2803 3418 2807
rect 3418 2803 3421 2807
rect 3342 2448 3346 2452
rect 3350 2428 3354 2432
rect 3310 2138 3314 2142
rect 3302 2078 3306 2082
rect 3294 2058 3298 2062
rect 3294 2048 3298 2052
rect 3302 1958 3306 1962
rect 3270 1878 3274 1882
rect 3270 1848 3274 1852
rect 3270 1798 3274 1802
rect 3326 2118 3330 2122
rect 3326 2068 3330 2072
rect 3358 2378 3362 2382
rect 3410 2603 3414 2607
rect 3417 2603 3418 2607
rect 3418 2603 3421 2607
rect 3414 2568 3418 2572
rect 3390 2478 3394 2482
rect 3398 2468 3402 2472
rect 3410 2403 3414 2407
rect 3417 2403 3418 2407
rect 3418 2403 3421 2407
rect 3494 2538 3498 2542
rect 3486 2468 3490 2472
rect 3430 2278 3434 2282
rect 3410 2203 3414 2207
rect 3417 2203 3418 2207
rect 3418 2203 3421 2207
rect 3374 2088 3378 2092
rect 3366 2078 3370 2082
rect 3350 2058 3354 2062
rect 3374 2058 3378 2062
rect 3230 1528 3234 1532
rect 3238 1488 3242 1492
rect 3262 1478 3266 1482
rect 3198 668 3202 672
rect 3182 558 3186 562
rect 3238 1168 3242 1172
rect 3238 1158 3242 1162
rect 3158 528 3162 532
rect 3182 278 3186 282
rect 3174 268 3178 272
rect 3158 148 3162 152
rect 3142 78 3146 82
rect 3270 1328 3274 1332
rect 3334 1858 3338 1862
rect 3318 1658 3322 1662
rect 3410 2003 3414 2007
rect 3417 2003 3418 2007
rect 3418 2003 3421 2007
rect 3390 1988 3394 1992
rect 3350 1528 3354 1532
rect 3294 1508 3298 1512
rect 3326 1508 3330 1512
rect 3414 1928 3418 1932
rect 3382 1838 3386 1842
rect 3398 1838 3402 1842
rect 3318 1378 3322 1382
rect 3374 1358 3378 1362
rect 3318 1348 3322 1352
rect 3262 928 3266 932
rect 3334 1288 3338 1292
rect 3358 1258 3362 1262
rect 3410 1803 3414 1807
rect 3417 1803 3418 1807
rect 3418 1803 3421 1807
rect 3438 2058 3442 2062
rect 3438 2018 3442 2022
rect 3446 1978 3450 1982
rect 3438 1928 3442 1932
rect 3430 1728 3434 1732
rect 3398 1688 3402 1692
rect 3398 1658 3402 1662
rect 3326 1148 3330 1152
rect 3390 1148 3394 1152
rect 3326 998 3330 1002
rect 3302 968 3306 972
rect 3382 1128 3386 1132
rect 3358 1058 3362 1062
rect 3350 1048 3354 1052
rect 3334 738 3338 742
rect 3294 718 3298 722
rect 3286 688 3290 692
rect 3278 498 3282 502
rect 3326 718 3330 722
rect 3310 598 3314 602
rect 3334 648 3338 652
rect 3318 408 3322 412
rect 3334 358 3338 362
rect 3294 158 3298 162
rect 3382 888 3386 892
rect 3382 718 3386 722
rect 3410 1603 3414 1607
rect 3417 1603 3418 1607
rect 3418 1603 3421 1607
rect 3462 2418 3466 2422
rect 3462 2288 3466 2292
rect 3462 2048 3466 2052
rect 3438 1468 3442 1472
rect 3454 1468 3458 1472
rect 3410 1403 3414 1407
rect 3417 1403 3418 1407
rect 3418 1403 3421 1407
rect 3422 1368 3426 1372
rect 3410 1203 3414 1207
rect 3417 1203 3418 1207
rect 3418 1203 3421 1207
rect 3430 1088 3434 1092
rect 3430 1068 3434 1072
rect 3410 1003 3414 1007
rect 3417 1003 3418 1007
rect 3418 1003 3421 1007
rect 3406 828 3410 832
rect 3410 803 3414 807
rect 3417 803 3418 807
rect 3418 803 3421 807
rect 3366 548 3370 552
rect 3366 528 3370 532
rect 3382 518 3386 522
rect 3366 148 3370 152
rect 3358 68 3362 72
rect 3410 603 3414 607
rect 3417 603 3418 607
rect 3418 603 3421 607
rect 3398 578 3402 582
rect 3430 558 3434 562
rect 3422 508 3426 512
rect 3454 1428 3458 1432
rect 3454 758 3458 762
rect 3446 748 3450 752
rect 3438 528 3442 532
rect 3410 403 3414 407
rect 3417 403 3418 407
rect 3418 403 3421 407
rect 3410 203 3414 207
rect 3417 203 3418 207
rect 3418 203 3421 207
rect 3414 138 3418 142
rect 3454 678 3458 682
rect 3462 528 3466 532
rect 3462 378 3466 382
rect 3486 2088 3490 2092
rect 3478 1888 3482 1892
rect 3486 1588 3490 1592
rect 3478 968 3482 972
rect 3478 818 3482 822
rect 3486 438 3490 442
rect 3518 2758 3522 2762
rect 3574 3478 3578 3482
rect 3510 2578 3514 2582
rect 3510 1958 3514 1962
rect 3574 2748 3578 2752
rect 3558 2648 3562 2652
rect 3566 2558 3570 2562
rect 3534 2118 3538 2122
rect 3526 2078 3530 2082
rect 3566 2308 3570 2312
rect 3558 2248 3562 2252
rect 3566 2138 3570 2142
rect 3542 1758 3546 1762
rect 3526 1718 3530 1722
rect 3534 1708 3538 1712
rect 3510 1558 3514 1562
rect 3510 1348 3514 1352
rect 3502 1338 3506 1342
rect 3510 1318 3514 1322
rect 3510 1078 3514 1082
rect 3510 858 3514 862
rect 3510 828 3514 832
rect 3510 548 3514 552
rect 3502 538 3506 542
rect 3510 498 3514 502
rect 3558 1928 3562 1932
rect 3566 1848 3570 1852
rect 3558 1838 3562 1842
rect 3574 1648 3578 1652
rect 3534 1468 3538 1472
rect 3542 1358 3546 1362
rect 3534 1138 3538 1142
rect 3590 3358 3594 3362
rect 3590 2758 3594 2762
rect 3590 2488 3594 2492
rect 3614 3088 3618 3092
rect 3622 3078 3626 3082
rect 3606 2148 3610 2152
rect 3606 2138 3610 2142
rect 3590 1658 3594 1662
rect 3590 1648 3594 1652
rect 3582 1368 3586 1372
rect 3574 1338 3578 1342
rect 3566 1258 3570 1262
rect 3582 1158 3586 1162
rect 3550 958 3554 962
rect 3518 418 3522 422
rect 3550 758 3554 762
rect 3542 748 3546 752
rect 3534 678 3538 682
rect 3558 628 3562 632
rect 3558 548 3562 552
rect 3558 528 3562 532
rect 3550 478 3554 482
rect 3550 348 3554 352
rect 3598 1488 3602 1492
rect 3622 2028 3626 2032
rect 3614 1938 3618 1942
rect 3622 1838 3626 1842
rect 3606 1438 3610 1442
rect 3622 1438 3626 1442
rect 3614 1388 3618 1392
rect 3606 1288 3610 1292
rect 3590 1118 3594 1122
rect 3582 708 3586 712
rect 3622 1258 3626 1262
rect 3606 1068 3610 1072
rect 3606 998 3610 1002
rect 3582 588 3586 592
rect 3590 328 3594 332
rect 3558 168 3562 172
rect 3574 168 3578 172
rect 3558 158 3562 162
rect 3622 988 3626 992
rect 3646 3438 3650 3442
rect 3646 3098 3650 3102
rect 3646 2748 3650 2752
rect 3654 2648 3658 2652
rect 3718 3528 3722 3532
rect 3670 3438 3674 3442
rect 3694 3368 3698 3372
rect 3710 3098 3714 3102
rect 3726 3088 3730 3092
rect 3702 3078 3706 3082
rect 3670 2418 3674 2422
rect 3694 2368 3698 2372
rect 3686 2278 3690 2282
rect 3702 2288 3706 2292
rect 3702 2278 3706 2282
rect 3670 2058 3674 2062
rect 3654 2048 3658 2052
rect 3646 1608 3650 1612
rect 3646 1368 3650 1372
rect 3654 1358 3658 1362
rect 3654 1348 3658 1352
rect 3654 1278 3658 1282
rect 3646 1158 3650 1162
rect 3630 888 3634 892
rect 3622 828 3626 832
rect 3614 748 3618 752
rect 3614 728 3618 732
rect 3614 708 3618 712
rect 3670 1508 3674 1512
rect 3686 1948 3690 1952
rect 3710 2138 3714 2142
rect 3710 1948 3714 1952
rect 3702 1728 3706 1732
rect 3686 1538 3690 1542
rect 3710 1568 3714 1572
rect 3678 1498 3682 1502
rect 3694 1488 3698 1492
rect 3702 1468 3706 1472
rect 3686 1438 3690 1442
rect 3686 1418 3690 1422
rect 3670 1338 3674 1342
rect 3670 1328 3674 1332
rect 3662 918 3666 922
rect 3654 888 3658 892
rect 3630 588 3634 592
rect 3638 508 3642 512
rect 3622 358 3626 362
rect 3630 358 3634 362
rect 3630 338 3634 342
rect 3622 248 3626 252
rect 3590 68 3594 72
rect 3478 58 3482 62
rect 3334 38 3338 42
rect 3390 38 3394 42
rect 3662 818 3666 822
rect 3654 508 3658 512
rect 3654 488 3658 492
rect 3654 448 3658 452
rect 3686 1268 3690 1272
rect 3686 1248 3690 1252
rect 3702 1438 3706 1442
rect 3670 648 3674 652
rect 3670 638 3674 642
rect 3670 368 3674 372
rect 3678 148 3682 152
rect 3742 3478 3746 3482
rect 3742 3448 3746 3452
rect 3734 2548 3738 2552
rect 3734 2028 3738 2032
rect 3734 1688 3738 1692
rect 3734 1598 3738 1602
rect 3726 1538 3730 1542
rect 3726 1418 3730 1422
rect 3726 1368 3730 1372
rect 3718 1318 3722 1322
rect 3710 658 3714 662
rect 3710 388 3714 392
rect 3710 348 3714 352
rect 3718 168 3722 172
rect 3718 158 3722 162
rect 3702 128 3706 132
rect 3718 78 3722 82
rect 3734 778 3738 782
rect 3734 768 3738 772
rect 3758 1948 3762 1952
rect 3758 1928 3762 1932
rect 3758 1858 3762 1862
rect 3750 1738 3754 1742
rect 3750 1638 3754 1642
rect 3758 1458 3762 1462
rect 3750 1248 3754 1252
rect 3758 1208 3762 1212
rect 3758 768 3762 772
rect 3750 338 3754 342
rect 3758 78 3762 82
rect 3774 1428 3778 1432
rect 346 3 350 7
rect 353 3 354 7
rect 354 3 357 7
rect 1362 3 1366 7
rect 1369 3 1370 7
rect 1370 3 1373 7
rect 2386 3 2390 7
rect 2393 3 2394 7
rect 2394 3 2397 7
rect 3410 3 3414 7
rect 3417 3 3418 7
rect 3418 3 3421 7
<< metal5 >>
rect 350 3603 353 3607
rect 349 3602 354 3603
rect 359 3602 360 3607
rect 1366 3603 1369 3607
rect 1365 3602 1370 3603
rect 1375 3602 1376 3607
rect 2390 3603 2393 3607
rect 2389 3602 2394 3603
rect 2399 3602 2400 3607
rect 3414 3603 3417 3607
rect 3413 3602 3418 3603
rect 3423 3602 3424 3607
rect 3570 3548 3606 3551
rect 914 3538 1390 3541
rect 2002 3538 2390 3541
rect 3218 3538 3318 3541
rect 3322 3538 3486 3541
rect 1806 3532 1809 3538
rect 3618 3538 3646 3541
rect 2274 3528 2574 3531
rect 3042 3528 3718 3531
rect 3722 3528 3741 3531
rect 1298 3518 1974 3521
rect 2242 3518 2494 3521
rect 3506 3518 3598 3521
rect 854 3503 857 3507
rect 853 3502 858 3503
rect 863 3502 864 3507
rect 1886 3503 1889 3507
rect 1885 3502 1890 3503
rect 1895 3502 1896 3507
rect 2910 3503 2913 3507
rect 2909 3502 2914 3503
rect 2919 3502 2920 3507
rect 986 3478 1870 3481
rect 3578 3478 3742 3481
rect 1170 3468 1414 3471
rect 2274 3458 2542 3461
rect 2578 3458 2958 3461
rect 2962 3458 3014 3461
rect 3742 3452 3745 3457
rect 2898 3448 3198 3451
rect 3602 3438 3646 3441
rect 3666 3438 3670 3441
rect 778 3418 2214 3421
rect 350 3403 353 3407
rect 349 3402 354 3403
rect 359 3402 360 3407
rect 1366 3403 1369 3407
rect 1365 3402 1370 3403
rect 1375 3402 1376 3407
rect 2390 3403 2393 3407
rect 2389 3402 2394 3403
rect 2399 3402 2400 3407
rect 3414 3403 3417 3407
rect 3413 3402 3418 3403
rect 3423 3402 3424 3407
rect 1562 3368 1646 3371
rect 3518 3361 3521 3368
rect 3274 3358 3521 3361
rect 3694 3361 3697 3368
rect 3594 3358 3697 3361
rect 1434 3348 1918 3351
rect 1122 3338 1350 3341
rect 3178 3338 3422 3341
rect 2130 3318 2294 3321
rect 2378 3308 2662 3311
rect 854 3303 857 3307
rect 853 3302 858 3303
rect 863 3302 864 3307
rect 1886 3303 1889 3307
rect 1885 3302 1890 3303
rect 1895 3302 1896 3307
rect 2910 3303 2913 3307
rect 2909 3302 2914 3303
rect 2919 3302 2920 3307
rect 1782 3281 1785 3288
rect 1186 3278 1785 3281
rect 146 3268 982 3271
rect 1298 3268 1646 3271
rect 1410 3258 1894 3261
rect 1298 3248 2966 3251
rect 2970 3248 3374 3251
rect 514 3238 2902 3241
rect 350 3203 353 3207
rect 349 3202 354 3203
rect 359 3202 360 3207
rect 1366 3203 1369 3207
rect 1365 3202 1370 3203
rect 1375 3202 1376 3207
rect 2390 3203 2393 3207
rect 2389 3202 2394 3203
rect 2399 3202 2400 3207
rect 3414 3203 3417 3207
rect 3413 3202 3418 3203
rect 3423 3202 3424 3207
rect 1002 3168 1798 3171
rect 978 3158 2222 3161
rect 3146 3158 3342 3161
rect 1554 3138 2294 3141
rect 2314 3138 2326 3141
rect 2202 3128 3118 3131
rect 1426 3118 2686 3121
rect 2234 3108 2470 3111
rect 854 3103 857 3107
rect 853 3102 858 3103
rect 863 3102 864 3107
rect 1886 3103 1889 3107
rect 1885 3102 1890 3103
rect 1895 3102 1896 3107
rect 2910 3103 2913 3107
rect 2909 3102 2914 3103
rect 2919 3102 2920 3107
rect 3646 3092 3649 3098
rect 3710 3092 3713 3098
rect 1738 3088 2126 3091
rect 3586 3088 3614 3091
rect 3726 3082 3729 3088
rect 2042 3078 2286 3081
rect 3626 3078 3693 3081
rect 3698 3078 3702 3081
rect 1998 3058 2078 3061
rect 2450 3058 2606 3061
rect 1042 3048 1230 3051
rect 1598 3051 1601 3058
rect 1998 3052 2001 3058
rect 1598 3048 1678 3051
rect 2066 3048 2166 3051
rect 2242 3048 2366 3051
rect 2370 3048 2462 3051
rect 898 3038 2270 3041
rect 2274 3038 2294 3041
rect 602 3028 2662 3031
rect 1802 3018 3030 3021
rect 1626 3008 2326 3011
rect 350 3003 353 3007
rect 349 3002 354 3003
rect 359 3002 360 3007
rect 1366 3003 1369 3007
rect 1365 3002 1370 3003
rect 1375 3002 1376 3007
rect 2390 3003 2393 3007
rect 2389 3002 2394 3003
rect 2399 3002 2400 3007
rect 3414 3003 3417 3007
rect 3413 3002 3418 3003
rect 3423 3002 3424 3007
rect 674 2988 950 2991
rect 1674 2988 2574 2991
rect 1554 2978 2014 2981
rect 2018 2978 2054 2981
rect 2058 2978 2118 2981
rect 2138 2978 3054 2981
rect 3194 2978 3470 2981
rect 1258 2968 1958 2971
rect 1962 2968 1974 2971
rect 2218 2968 2310 2971
rect 3122 2968 3502 2971
rect 1226 2958 1289 2961
rect 1322 2958 1654 2961
rect 1666 2958 2822 2961
rect 1286 2952 1289 2958
rect 1730 2948 2270 2951
rect 3330 2948 3374 2951
rect 754 2938 1246 2941
rect 1594 2938 1846 2941
rect 2130 2938 2318 2941
rect 2378 2938 2702 2941
rect 1634 2928 2006 2931
rect 2010 2928 2209 2931
rect 2342 2928 2350 2931
rect 2354 2928 2502 2931
rect 2206 2922 2209 2928
rect 1306 2918 1702 2921
rect 1842 2918 1902 2921
rect 2138 2908 2350 2911
rect 854 2903 857 2907
rect 853 2902 858 2903
rect 863 2902 864 2907
rect 1886 2903 1889 2907
rect 1885 2902 1890 2903
rect 1895 2902 1896 2907
rect 2910 2903 2913 2907
rect 2909 2902 2914 2903
rect 2919 2902 2920 2907
rect 1506 2888 2582 2891
rect 1478 2881 1481 2888
rect 1478 2878 2054 2881
rect 2266 2878 2790 2881
rect 770 2868 790 2871
rect 794 2868 854 2871
rect 1498 2868 2070 2871
rect 2074 2868 2390 2871
rect 2458 2868 2694 2871
rect 770 2858 1302 2861
rect 2074 2858 2158 2861
rect 42 2848 118 2851
rect 258 2848 1118 2851
rect 2662 2851 2665 2858
rect 2338 2848 2665 2851
rect 1866 2828 2550 2831
rect 1186 2818 1766 2821
rect 1770 2818 3414 2821
rect 350 2803 353 2807
rect 349 2802 354 2803
rect 359 2802 360 2807
rect 1366 2803 1369 2807
rect 1365 2802 1370 2803
rect 1375 2802 1376 2807
rect 1790 2802 1793 2808
rect 2390 2803 2393 2807
rect 2389 2802 2394 2803
rect 2399 2802 2400 2807
rect 3414 2803 3417 2807
rect 3413 2802 3418 2803
rect 3423 2802 3424 2807
rect 1490 2798 1670 2801
rect 1794 2798 2350 2801
rect 818 2788 990 2791
rect 1130 2788 2918 2791
rect 834 2778 894 2781
rect 1714 2778 1982 2781
rect 762 2768 806 2771
rect 1018 2768 1734 2771
rect 1746 2768 1990 2771
rect 1018 2758 1150 2761
rect 1618 2758 1870 2761
rect 3026 2758 3518 2761
rect 3522 2758 3590 2761
rect 138 2748 1702 2751
rect 1738 2748 2030 2751
rect 3458 2748 3574 2751
rect 3578 2748 3646 2751
rect 1666 2738 1814 2741
rect 878 2731 881 2738
rect 826 2728 881 2731
rect 1594 2728 1742 2731
rect 1810 2728 1814 2731
rect 842 2718 894 2721
rect 1650 2718 2446 2721
rect 2866 2718 3270 2721
rect 1946 2708 2454 2711
rect 2458 2708 2766 2711
rect 854 2703 857 2707
rect 853 2702 858 2703
rect 863 2702 864 2707
rect 1886 2703 1889 2707
rect 1885 2702 1890 2703
rect 1895 2702 1896 2707
rect 2910 2703 2913 2707
rect 2909 2702 2914 2703
rect 2919 2702 2920 2707
rect 946 2698 1830 2701
rect 802 2688 974 2691
rect 1874 2688 2270 2691
rect 2274 2688 2822 2691
rect 758 2678 766 2681
rect 1086 2681 1089 2688
rect 770 2678 1089 2681
rect 1826 2678 1958 2681
rect 2402 2678 3110 2681
rect 506 2668 878 2671
rect 1706 2668 2150 2671
rect 2410 2668 2902 2671
rect 730 2658 1030 2661
rect 2114 2658 3174 2661
rect 674 2648 881 2651
rect 1794 2648 2414 2651
rect 2690 2648 2774 2651
rect 2834 2648 2894 2651
rect 3562 2648 3654 2651
rect 878 2642 881 2648
rect 378 2638 726 2641
rect 1930 2638 2686 2641
rect 2690 2638 2758 2641
rect 482 2628 798 2631
rect 858 2628 1006 2631
rect 2130 2618 2926 2621
rect 1698 2608 1886 2611
rect 350 2603 353 2607
rect 349 2602 354 2603
rect 359 2602 360 2607
rect 1366 2603 1369 2607
rect 1365 2602 1370 2603
rect 1375 2602 1376 2607
rect 2390 2603 2393 2607
rect 2389 2602 2394 2603
rect 2399 2602 2400 2607
rect 3414 2603 3417 2607
rect 3413 2602 3418 2603
rect 3423 2602 3424 2607
rect 2650 2598 3262 2601
rect 2522 2578 2998 2581
rect 3002 2578 3510 2581
rect 2770 2568 2790 2571
rect 2802 2568 3150 2571
rect 3154 2568 3414 2571
rect 646 2561 649 2568
rect 646 2558 662 2561
rect 1026 2558 1630 2561
rect 1830 2558 2062 2561
rect 2466 2558 3102 2561
rect 3242 2558 3566 2561
rect 1830 2552 1833 2558
rect 802 2548 910 2551
rect 1762 2548 1814 2551
rect 2410 2548 2510 2551
rect 878 2538 1094 2541
rect 1730 2538 1854 2541
rect 1858 2538 2590 2541
rect 878 2532 881 2538
rect 3186 2538 3494 2541
rect 3734 2541 3737 2548
rect 3730 2538 3737 2541
rect 1626 2528 2238 2531
rect 2298 2528 3070 2531
rect 2442 2518 2814 2521
rect 854 2503 857 2507
rect 853 2502 858 2503
rect 863 2502 864 2507
rect 1886 2503 1889 2507
rect 1885 2502 1890 2503
rect 1895 2502 1896 2507
rect 2910 2503 2913 2507
rect 2909 2502 2914 2503
rect 2919 2502 2920 2507
rect 1914 2498 2366 2501
rect 138 2488 982 2491
rect 1786 2488 1910 2491
rect 1914 2488 2414 2491
rect 3122 2488 3230 2491
rect 3258 2488 3590 2491
rect 2546 2478 2862 2481
rect 3074 2478 3390 2481
rect 546 2468 734 2471
rect 842 2468 1214 2471
rect 3402 2468 3486 2471
rect 994 2458 1137 2461
rect 1134 2452 1137 2458
rect 1198 2458 1566 2461
rect 1198 2452 1201 2458
rect 2154 2448 2990 2451
rect 3274 2448 3342 2451
rect 194 2438 1214 2441
rect 1242 2428 3350 2431
rect 3122 2418 3462 2421
rect 3474 2418 3670 2421
rect 350 2403 353 2407
rect 349 2402 354 2403
rect 359 2402 360 2407
rect 1366 2403 1369 2407
rect 1365 2402 1370 2403
rect 1375 2402 1376 2407
rect 2390 2403 2393 2407
rect 2389 2402 2394 2403
rect 2399 2402 2400 2407
rect 3414 2403 3417 2407
rect 3413 2402 3418 2403
rect 3423 2402 3424 2407
rect 1970 2388 3270 2391
rect 1722 2378 2598 2381
rect 2714 2378 3358 2381
rect 650 2368 678 2371
rect 1842 2368 2166 2371
rect 2642 2368 3118 2371
rect 3634 2368 3694 2371
rect 1242 2358 1598 2361
rect 1002 2348 1294 2351
rect 1434 2348 2526 2351
rect 1490 2338 1854 2341
rect 2322 2338 2406 2341
rect 2626 2338 2830 2341
rect 2998 2341 3001 2348
rect 2858 2338 3001 2341
rect 1234 2328 2806 2331
rect 2810 2328 2870 2331
rect 1722 2318 2030 2321
rect 2338 2318 2470 2321
rect 2866 2318 2926 2321
rect 2146 2308 2606 2311
rect 3226 2308 3566 2311
rect 854 2303 857 2307
rect 853 2302 858 2303
rect 863 2302 864 2307
rect 1886 2303 1889 2307
rect 1885 2302 1890 2303
rect 1895 2302 1896 2307
rect 2910 2303 2913 2307
rect 2909 2302 2914 2303
rect 2919 2302 2920 2307
rect 2010 2298 2893 2301
rect 1738 2288 3054 2291
rect 3058 2288 3462 2291
rect 3682 2288 3702 2291
rect 1450 2278 1485 2281
rect 1554 2278 2254 2281
rect 2258 2278 2438 2281
rect 3170 2278 3430 2281
rect 3462 2278 3686 2281
rect 1502 2271 1505 2278
rect 1098 2268 1505 2271
rect 1514 2268 1782 2271
rect 1850 2268 2182 2271
rect 2186 2268 2310 2271
rect 2490 2268 2622 2271
rect 3462 2271 3465 2278
rect 3698 2278 3702 2281
rect 2898 2268 3465 2271
rect 3206 2262 3209 2268
rect 1362 2258 1990 2261
rect 1994 2258 2150 2261
rect 2378 2258 2550 2261
rect 2554 2258 3038 2261
rect 762 2248 1078 2251
rect 1858 2248 2478 2251
rect 3522 2248 3558 2251
rect 1314 2228 2014 2231
rect 1562 2218 3270 2221
rect 1770 2208 2022 2211
rect 2026 2208 2230 2211
rect 2234 2208 2358 2211
rect 350 2203 353 2207
rect 349 2202 354 2203
rect 359 2202 360 2207
rect 1366 2203 1369 2207
rect 1365 2202 1370 2203
rect 1375 2202 1376 2207
rect 2390 2203 2393 2207
rect 2389 2202 2394 2203
rect 2399 2202 2400 2207
rect 3414 2203 3417 2207
rect 3413 2202 3418 2203
rect 3423 2202 3424 2207
rect 1738 2188 2022 2191
rect 1450 2178 1702 2181
rect 1706 2178 1846 2181
rect 1850 2178 1902 2181
rect 2154 2178 3110 2181
rect 1130 2168 1390 2171
rect 1514 2168 2510 2171
rect 1162 2158 2094 2161
rect 2450 2158 2534 2161
rect 1858 2148 1926 2151
rect 2098 2148 2942 2151
rect 3610 2148 3713 2151
rect 3710 2142 3713 2148
rect 134 2138 750 2141
rect 970 2138 1614 2141
rect 2786 2138 2822 2141
rect 3314 2138 3566 2141
rect 3610 2138 3661 2141
rect 134 2132 137 2138
rect 2874 2128 2966 2131
rect 2210 2118 2766 2121
rect 2826 2118 3326 2121
rect 3330 2118 3534 2121
rect 854 2103 857 2107
rect 853 2102 858 2103
rect 863 2102 864 2107
rect 1886 2103 1889 2107
rect 1885 2102 1890 2103
rect 1895 2102 1896 2107
rect 2910 2103 2913 2107
rect 2909 2102 2914 2103
rect 2919 2102 2920 2107
rect 2546 2098 2806 2101
rect 1178 2088 2590 2091
rect 2610 2088 3078 2091
rect 3378 2088 3486 2091
rect 2434 2078 2582 2081
rect 3306 2078 3366 2081
rect 3530 2078 3533 2081
rect 1738 2068 2182 2071
rect 2234 2068 3326 2071
rect 1154 2058 1438 2061
rect 1938 2058 2526 2061
rect 2594 2058 2830 2061
rect 3298 2058 3350 2061
rect 3378 2058 3438 2061
rect 3666 2058 3670 2061
rect 1794 2048 1801 2051
rect 2210 2048 2494 2051
rect 3298 2048 3462 2051
rect 1798 2042 1801 2048
rect 2290 2038 2670 2041
rect 3654 2041 3657 2048
rect 3698 2048 3709 2051
rect 2690 2038 3657 2041
rect 3714 2038 3737 2041
rect 3734 2032 3737 2038
rect 1834 2028 2854 2031
rect 3442 2028 3622 2031
rect 1842 2018 3438 2021
rect 2410 2008 2846 2011
rect 350 2003 353 2007
rect 349 2002 354 2003
rect 359 2002 360 2007
rect 1366 2003 1369 2007
rect 1365 2002 1370 2003
rect 1375 2002 1376 2007
rect 2390 2003 2393 2007
rect 2389 2002 2394 2003
rect 2399 2002 2400 2007
rect 3414 2003 3417 2007
rect 3413 2002 3418 2003
rect 3423 2002 3424 2007
rect 2322 1988 3390 1991
rect 1930 1978 3166 1981
rect 3170 1978 3446 1981
rect 2802 1968 2934 1971
rect 10 1958 990 1961
rect 2378 1958 3302 1961
rect 3306 1958 3510 1961
rect 50 1948 734 1951
rect 842 1948 998 1951
rect 1282 1948 2462 1951
rect 2746 1948 3006 1951
rect 3074 1948 3161 1951
rect 3158 1942 3161 1948
rect 3618 1948 3686 1951
rect 3714 1948 3758 1951
rect 202 1938 478 1941
rect 714 1938 758 1941
rect 1570 1938 1686 1941
rect 1778 1938 2310 1941
rect 3130 1938 3133 1941
rect 3614 1932 3617 1938
rect 3758 1932 3761 1937
rect 1586 1928 1630 1931
rect 2762 1928 2958 1931
rect 2962 1928 3414 1931
rect 3442 1928 3558 1931
rect 1810 1918 2126 1921
rect 2890 1918 3054 1921
rect 854 1903 857 1907
rect 853 1902 858 1903
rect 863 1902 864 1907
rect 1886 1903 1889 1907
rect 1885 1902 1890 1903
rect 1895 1902 1896 1907
rect 2910 1903 2913 1907
rect 2909 1902 2914 1903
rect 2919 1902 2920 1907
rect 1474 1898 1598 1901
rect 786 1888 1430 1891
rect 2178 1888 2438 1891
rect 1202 1878 1510 1881
rect 2034 1878 2198 1881
rect 2282 1878 2302 1881
rect 2346 1878 2454 1881
rect 3478 1881 3481 1888
rect 3274 1878 3481 1881
rect 1674 1868 2374 1871
rect 2922 1868 2998 1871
rect 3758 1868 3773 1871
rect 3758 1862 3761 1868
rect 2354 1858 2534 1861
rect 2538 1858 2654 1861
rect 3106 1858 3334 1861
rect 18 1848 606 1851
rect 610 1848 918 1851
rect 1962 1848 2414 1851
rect 2458 1848 2758 1851
rect 3274 1848 3566 1851
rect 1594 1838 3150 1841
rect 3154 1838 3382 1841
rect 3402 1838 3558 1841
rect 3570 1838 3622 1841
rect 2814 1822 2817 1828
rect 1794 1818 2630 1821
rect 2682 1808 2702 1811
rect 350 1803 353 1807
rect 349 1802 354 1803
rect 359 1802 360 1807
rect 1366 1803 1369 1807
rect 1365 1802 1370 1803
rect 1375 1802 1376 1807
rect 2390 1803 2393 1807
rect 2389 1802 2394 1803
rect 2399 1802 2400 1807
rect 3414 1803 3417 1807
rect 3413 1802 3418 1803
rect 3423 1802 3424 1807
rect 1682 1798 2070 1801
rect 2074 1798 2377 1801
rect 3242 1798 3270 1801
rect 2010 1788 2318 1791
rect 2374 1791 2377 1798
rect 2374 1788 2710 1791
rect 2274 1778 3126 1781
rect 1578 1768 3158 1771
rect 1378 1758 2374 1761
rect 2394 1758 2758 1761
rect 3546 1758 3581 1761
rect 2370 1748 2750 1751
rect 2862 1751 2865 1758
rect 2862 1748 2982 1751
rect 3378 1748 3753 1751
rect 3750 1742 3753 1748
rect 482 1738 654 1741
rect 658 1738 814 1741
rect 1338 1738 1638 1741
rect 2674 1738 2710 1741
rect 2714 1738 2870 1741
rect 138 1728 1054 1731
rect 1874 1728 1993 1731
rect 2138 1728 3230 1731
rect 3242 1728 3430 1731
rect 3706 1728 3725 1731
rect 1990 1722 1993 1728
rect 778 1718 926 1721
rect 946 1718 1926 1721
rect 2402 1718 3526 1721
rect 3162 1708 3534 1711
rect 854 1703 857 1707
rect 853 1702 858 1703
rect 863 1702 864 1707
rect 1886 1703 1889 1707
rect 1885 1702 1890 1703
rect 1895 1702 1896 1707
rect 2910 1703 2913 1707
rect 2909 1702 2914 1703
rect 2919 1702 2920 1707
rect 914 1688 1054 1691
rect 2050 1688 2366 1691
rect 2850 1688 2990 1691
rect 3006 1688 3398 1691
rect 3006 1681 3009 1688
rect 3554 1688 3734 1691
rect 1914 1678 3009 1681
rect 122 1668 998 1671
rect 1038 1671 1041 1678
rect 1038 1668 1350 1671
rect 2778 1668 2838 1671
rect 3010 1668 3086 1671
rect 10 1658 526 1661
rect 1098 1658 1494 1661
rect 2650 1658 3318 1661
rect 3402 1658 3590 1661
rect 946 1648 1326 1651
rect 3578 1648 3590 1651
rect 986 1638 1206 1641
rect 3714 1638 3750 1641
rect 98 1628 1638 1631
rect 1026 1618 1614 1621
rect 3570 1608 3646 1611
rect 350 1603 353 1607
rect 349 1602 354 1603
rect 359 1602 360 1607
rect 1366 1603 1369 1607
rect 1365 1602 1370 1603
rect 1375 1602 1376 1607
rect 2390 1603 2393 1607
rect 2389 1602 2394 1603
rect 2399 1602 2400 1607
rect 3414 1603 3417 1607
rect 3413 1602 3418 1603
rect 3423 1602 3424 1607
rect 3738 1598 3741 1601
rect 3074 1588 3190 1591
rect 3194 1588 3486 1591
rect 3130 1568 3133 1571
rect 1186 1558 1958 1561
rect 3126 1561 3129 1568
rect 3710 1562 3713 1568
rect 2810 1558 3129 1561
rect 1074 1548 1406 1551
rect 1410 1548 1581 1551
rect 1586 1548 1606 1551
rect 3510 1551 3513 1558
rect 3510 1548 3533 1551
rect 3506 1538 3533 1541
rect 3690 1538 3726 1541
rect 3234 1528 3350 1531
rect 834 1518 3070 1521
rect 2698 1508 2854 1511
rect 3298 1508 3326 1511
rect 3674 1508 3677 1511
rect 854 1503 857 1507
rect 853 1502 858 1503
rect 863 1502 864 1507
rect 1886 1503 1889 1507
rect 1885 1502 1890 1503
rect 1895 1502 1896 1507
rect 2910 1503 2913 1507
rect 2909 1502 2914 1503
rect 2919 1502 2920 1507
rect 2714 1498 2870 1501
rect 3678 1492 3681 1498
rect 1946 1488 2590 1491
rect 2610 1488 3238 1491
rect 3490 1488 3598 1491
rect 3694 1482 3697 1488
rect 1330 1478 1878 1481
rect 1882 1478 2486 1481
rect 2594 1478 3110 1481
rect 3170 1478 3262 1481
rect 666 1468 974 1471
rect 978 1468 1062 1471
rect 2858 1468 3006 1471
rect 3442 1468 3454 1471
rect 3538 1468 3702 1471
rect 1058 1458 1550 1461
rect 3634 1458 3758 1461
rect 1042 1448 1910 1451
rect 2058 1448 2758 1451
rect 3602 1448 3629 1451
rect 1634 1438 1942 1441
rect 3610 1438 3622 1441
rect 3690 1438 3702 1441
rect 1722 1428 3062 1431
rect 3458 1428 3774 1431
rect 1682 1418 3206 1421
rect 3690 1418 3726 1421
rect 1386 1408 1886 1411
rect 350 1403 353 1407
rect 349 1402 354 1403
rect 359 1402 360 1407
rect 1366 1403 1369 1407
rect 1365 1402 1370 1403
rect 1375 1402 1376 1407
rect 2390 1403 2393 1407
rect 2389 1402 2394 1403
rect 2399 1402 2400 1407
rect 3414 1403 3417 1407
rect 3413 1402 3418 1403
rect 3423 1402 3424 1407
rect 666 1388 782 1391
rect 786 1388 1158 1391
rect 1306 1388 2166 1391
rect 2170 1388 2502 1391
rect 2506 1388 2958 1391
rect 3330 1388 3614 1391
rect 1618 1378 3318 1381
rect 3602 1378 3645 1381
rect 1706 1368 2566 1371
rect 2850 1368 3422 1371
rect 3586 1368 3646 1371
rect 1454 1361 1457 1368
rect 3698 1368 3726 1371
rect 538 1358 1870 1361
rect 1890 1358 2094 1361
rect 2274 1358 3374 1361
rect 3378 1358 3542 1361
rect 3650 1358 3654 1361
rect 1442 1348 1462 1351
rect 2066 1348 3318 1351
rect 3514 1348 3654 1351
rect 18 1338 558 1341
rect 1070 1341 1073 1348
rect 1070 1338 1270 1341
rect 1410 1338 2281 1341
rect 2278 1332 2281 1338
rect 3578 1338 3670 1341
rect 3502 1332 3505 1338
rect 482 1328 814 1331
rect 818 1328 1238 1331
rect 2490 1328 2798 1331
rect 2962 1328 3134 1331
rect 3138 1328 3270 1331
rect 3674 1328 3725 1331
rect 178 1318 1062 1321
rect 1842 1318 2326 1321
rect 2514 1318 3510 1321
rect 3634 1318 3718 1321
rect 970 1308 1622 1311
rect 2002 1308 2678 1311
rect 3154 1308 3174 1311
rect 854 1303 857 1307
rect 853 1302 858 1303
rect 863 1302 864 1307
rect 1886 1303 1889 1307
rect 1885 1302 1890 1303
rect 1895 1302 1896 1307
rect 2910 1303 2913 1307
rect 2909 1302 2914 1303
rect 2919 1302 2920 1307
rect 1346 1298 1838 1301
rect 2994 1298 3142 1301
rect 1266 1288 2294 1291
rect 2834 1288 2934 1291
rect 2938 1288 3334 1291
rect 3338 1288 3606 1291
rect 3066 1278 3069 1281
rect 3650 1278 3654 1281
rect 1954 1268 2342 1271
rect 3182 1268 3533 1271
rect 3182 1261 3185 1268
rect 3538 1268 3686 1271
rect 1666 1258 3185 1261
rect 3362 1258 3566 1261
rect 3626 1258 3645 1261
rect 1154 1248 2318 1251
rect 3186 1248 3686 1251
rect 3754 1248 3757 1251
rect 1410 1228 2982 1231
rect 3006 1222 3009 1228
rect 1170 1218 2646 1221
rect 350 1203 353 1207
rect 349 1202 354 1203
rect 359 1202 360 1207
rect 1366 1203 1369 1207
rect 1365 1202 1370 1203
rect 1375 1202 1376 1207
rect 2390 1203 2393 1207
rect 2389 1202 2394 1203
rect 2399 1202 2400 1207
rect 3414 1203 3417 1207
rect 3413 1202 3418 1203
rect 3423 1202 3424 1207
rect 3758 1202 3761 1208
rect 2426 1198 2950 1201
rect 1626 1188 1966 1191
rect 2578 1188 2966 1191
rect 1402 1178 1702 1181
rect 1738 1178 2374 1181
rect 2434 1178 2662 1181
rect 18 1168 558 1171
rect 1730 1168 2150 1171
rect 2482 1168 3238 1171
rect 2170 1158 2494 1161
rect 2498 1158 2638 1161
rect 3242 1158 3453 1161
rect 3586 1158 3646 1161
rect 18 1148 998 1151
rect 1442 1148 1801 1151
rect 2034 1148 3326 1151
rect 538 1138 702 1141
rect 1090 1138 1646 1141
rect 1798 1141 1801 1148
rect 3390 1142 3393 1148
rect 3534 1142 3537 1147
rect 1798 1138 2454 1141
rect 2490 1138 2934 1141
rect 1202 1128 1526 1131
rect 2218 1128 2550 1131
rect 2810 1128 3382 1131
rect 1266 1118 1470 1121
rect 1606 1118 2110 1121
rect 2442 1118 2518 1121
rect 3090 1118 3110 1121
rect 1606 1111 1609 1118
rect 3586 1118 3590 1121
rect 1250 1108 1609 1111
rect 1618 1108 1670 1111
rect 2042 1108 2126 1111
rect 2306 1108 2470 1111
rect 854 1103 857 1107
rect 853 1102 858 1103
rect 863 1102 864 1107
rect 1886 1103 1889 1107
rect 1885 1102 1890 1103
rect 1895 1102 1896 1107
rect 2910 1103 2913 1107
rect 2909 1102 2914 1103
rect 2919 1102 2920 1107
rect 3038 1102 3041 1108
rect 2058 1098 2478 1101
rect 1026 1088 1222 1091
rect 1226 1088 1438 1091
rect 2090 1088 3430 1091
rect 1114 1078 1230 1081
rect 1662 1078 1846 1081
rect 2186 1078 3510 1081
rect 1662 1072 1665 1078
rect 26 1068 894 1071
rect 938 1068 1350 1071
rect 1354 1068 1462 1071
rect 1602 1068 1638 1071
rect 2298 1068 2470 1071
rect 2602 1068 2806 1071
rect 2994 1068 3430 1071
rect 3610 1068 3773 1071
rect 58 1058 326 1061
rect 954 1058 990 1061
rect 1506 1058 1662 1061
rect 2186 1058 2598 1061
rect 3018 1058 3358 1061
rect 1098 1048 1350 1051
rect 1418 1048 2446 1051
rect 2450 1048 2566 1051
rect 2578 1048 2702 1051
rect 2762 1048 3038 1051
rect 3354 1048 3373 1051
rect 1162 1038 1638 1041
rect 2378 1038 2790 1041
rect 2866 1038 2982 1041
rect 2986 1038 3134 1041
rect 1162 1028 1830 1031
rect 1994 1028 2558 1031
rect 2562 1028 2958 1031
rect 1290 1018 1526 1021
rect 1530 1018 1766 1021
rect 1862 1018 3158 1021
rect 1862 1011 1865 1018
rect 1426 1008 1865 1011
rect 1874 1008 2166 1011
rect 3034 1008 3038 1011
rect 350 1003 353 1007
rect 349 1002 354 1003
rect 359 1002 360 1007
rect 1366 1003 1369 1007
rect 1365 1002 1370 1003
rect 1375 1002 1376 1007
rect 2390 1003 2393 1007
rect 2389 1002 2394 1003
rect 2399 1002 2400 1007
rect 3414 1003 3417 1007
rect 3413 1002 3418 1003
rect 3423 1002 3424 1007
rect 1554 998 1662 1001
rect 2146 998 2374 1001
rect 2498 998 2574 1001
rect 2646 998 3326 1001
rect 3610 998 3613 1001
rect 2646 991 2649 998
rect 1818 988 2649 991
rect 2666 988 2798 991
rect 2810 988 3118 991
rect 3618 988 3622 991
rect 2130 978 3134 981
rect 2578 968 3302 971
rect 1138 958 1726 961
rect 1962 958 2630 961
rect 2746 958 2974 961
rect 3478 961 3481 968
rect 3478 958 3550 961
rect 1490 948 1830 951
rect 1834 948 1870 951
rect 1874 948 2758 951
rect 2834 948 2862 951
rect 3062 951 3065 958
rect 2882 948 3065 951
rect 1858 938 1974 941
rect 2066 938 2286 941
rect 2066 928 2206 931
rect 2370 928 2877 931
rect 3074 928 3262 931
rect 1210 918 1958 921
rect 2642 918 3006 921
rect 3634 918 3662 921
rect 854 903 857 907
rect 853 902 858 903
rect 863 902 864 907
rect 1886 903 1889 907
rect 1885 902 1890 903
rect 1895 902 1896 907
rect 2910 903 2913 907
rect 2909 902 2914 903
rect 2919 902 2920 907
rect 322 898 542 901
rect 2194 898 2366 901
rect 2370 898 2598 901
rect 2770 888 3382 891
rect 3634 888 3654 891
rect 86 881 89 888
rect 86 878 566 881
rect 1898 878 2750 881
rect 2850 878 3006 881
rect 1034 868 1318 871
rect 1502 871 1505 878
rect 1502 868 1774 871
rect 2066 868 2510 871
rect 2714 868 2902 871
rect 2906 868 2942 871
rect 3006 871 3009 878
rect 3006 868 3150 871
rect 2586 858 2678 861
rect 2874 858 2918 861
rect 3074 858 3510 861
rect 1578 848 1822 851
rect 1930 848 2262 851
rect 2634 848 2854 851
rect 1490 838 2038 841
rect 1730 828 2478 831
rect 2482 828 2686 831
rect 2690 828 2822 831
rect 2842 828 3406 831
rect 3514 828 3622 831
rect 1818 818 2102 821
rect 2130 818 3478 821
rect 3482 818 3662 821
rect 1706 808 2214 811
rect 2906 808 2982 811
rect 350 803 353 807
rect 349 802 354 803
rect 359 802 360 807
rect 1366 803 1369 807
rect 1365 802 1370 803
rect 1375 802 1376 807
rect 2390 803 2393 807
rect 2389 802 2394 803
rect 2399 802 2400 807
rect 3414 803 3417 807
rect 3413 802 3418 803
rect 3423 802 3424 807
rect 1410 798 1862 801
rect 2434 798 2654 801
rect 1386 788 2134 791
rect 2218 788 2494 791
rect 1858 778 3022 781
rect 3730 778 3734 781
rect 1578 768 1646 771
rect 1650 768 1870 771
rect 2290 768 2518 771
rect 2754 768 3126 771
rect 3738 768 3758 771
rect 1602 758 2062 761
rect 3458 758 3550 761
rect 1510 751 1513 758
rect 1510 748 1558 751
rect 2258 748 2486 751
rect 2506 748 2678 751
rect 2698 748 2902 751
rect 3442 748 3446 751
rect 3546 748 3614 751
rect 1546 738 1918 741
rect 1938 738 3334 741
rect 3614 732 3617 737
rect 66 728 102 731
rect 2106 728 2518 731
rect 2858 728 2942 731
rect 2986 728 3086 731
rect 3090 728 3102 731
rect 826 718 2350 721
rect 2386 718 3294 721
rect 3330 718 3382 721
rect 3586 708 3614 711
rect 854 703 857 707
rect 853 702 858 703
rect 863 702 864 707
rect 1886 703 1889 707
rect 1885 702 1890 703
rect 1895 702 1896 707
rect 2910 703 2913 707
rect 2909 702 2914 703
rect 2919 702 2920 707
rect 3166 702 3169 708
rect 1914 698 2446 701
rect 2954 698 2966 701
rect 178 688 494 691
rect 1866 688 3286 691
rect 86 681 89 688
rect 3534 682 3537 687
rect 86 678 654 681
rect 1810 678 2022 681
rect 2026 678 2254 681
rect 2274 678 3454 681
rect 1602 668 1606 671
rect 2970 668 3198 671
rect 1926 661 1929 668
rect 1926 658 1958 661
rect 2106 658 2334 661
rect 3098 658 3149 661
rect 3154 658 3158 661
rect 3670 658 3710 661
rect 3670 652 3673 658
rect 1242 648 2102 651
rect 2234 648 2310 651
rect 2314 648 2486 651
rect 2778 648 3334 651
rect 2066 638 2414 641
rect 2706 638 2854 641
rect 3650 638 3670 641
rect 2090 628 3558 631
rect 2242 618 2526 621
rect 2530 618 2894 621
rect 2626 608 2806 611
rect 2850 608 3006 611
rect 350 603 353 607
rect 349 602 354 603
rect 359 602 360 607
rect 1366 603 1369 607
rect 1365 602 1370 603
rect 1375 602 1376 607
rect 2390 603 2393 607
rect 2389 602 2394 603
rect 2399 602 2400 607
rect 3414 603 3417 607
rect 3413 602 3418 603
rect 3423 602 3424 607
rect 1538 598 2374 601
rect 2522 598 2774 601
rect 2826 598 2950 601
rect 3130 598 3310 601
rect 1650 588 3118 591
rect 3586 588 3630 591
rect 1490 578 2742 581
rect 2746 578 2749 581
rect 2770 578 2998 581
rect 3182 578 3398 581
rect 1370 568 2038 571
rect 2042 568 2086 571
rect 3182 571 3185 578
rect 2162 568 3185 571
rect 2258 558 2686 561
rect 2778 558 2910 561
rect 3186 558 3430 561
rect 1330 548 1542 551
rect 1546 548 1581 551
rect 1594 548 1790 551
rect 1794 548 2078 551
rect 2082 548 2182 551
rect 2450 548 3366 551
rect 3514 548 3558 551
rect 914 538 1550 541
rect 2138 538 2334 541
rect 2722 538 2798 541
rect 2866 538 3070 541
rect 3074 538 3502 541
rect 2370 528 3158 531
rect 3370 528 3438 531
rect 3466 528 3558 531
rect 1434 518 2822 521
rect 2898 518 3382 521
rect 3114 508 3422 511
rect 3642 508 3654 511
rect 854 503 857 507
rect 853 502 858 503
rect 863 502 864 507
rect 1886 503 1889 507
rect 1885 502 1890 503
rect 1895 502 1896 507
rect 2910 503 2913 507
rect 2909 502 2914 503
rect 2919 502 2920 507
rect 3070 502 3073 507
rect 3282 498 3510 501
rect 386 488 790 491
rect 810 488 1606 491
rect 1610 488 1902 491
rect 2546 488 3654 491
rect 1866 478 3550 481
rect 1290 468 1510 471
rect 1834 468 1942 471
rect 2450 468 3110 471
rect 1258 458 1486 461
rect 2018 458 2254 461
rect 2370 458 2734 461
rect 2818 458 2822 461
rect 2858 458 2926 461
rect 2338 448 2462 451
rect 2754 448 3654 451
rect 2178 438 2382 441
rect 2494 438 2630 441
rect 2858 438 3486 441
rect 2494 431 2497 438
rect 1978 428 2497 431
rect 2790 431 2793 438
rect 2506 428 2793 431
rect 3518 422 3521 427
rect 1770 418 2878 421
rect 2466 408 3318 411
rect 350 403 353 407
rect 349 402 354 403
rect 359 402 360 407
rect 1366 403 1369 407
rect 1365 402 1370 403
rect 1375 402 1376 407
rect 2390 403 2393 407
rect 2389 402 2394 403
rect 2399 402 2400 407
rect 3414 403 3417 407
rect 3413 402 3418 403
rect 3423 402 3424 407
rect 1234 388 2046 391
rect 2210 388 3710 391
rect 1874 378 2782 381
rect 2786 378 3462 381
rect 1026 368 1102 371
rect 2018 368 2513 371
rect 2570 368 2862 371
rect 2510 362 2513 368
rect 3630 362 3633 367
rect 3338 358 3622 361
rect 3670 361 3673 368
rect 3666 358 3673 361
rect 1074 348 1942 351
rect 2034 348 2646 351
rect 2650 348 2718 351
rect 2754 348 2918 351
rect 3506 348 3550 351
rect 3602 348 3710 351
rect 546 338 934 341
rect 1554 338 1846 341
rect 2282 338 2326 341
rect 2354 338 2374 341
rect 3586 338 3630 341
rect 3634 338 3750 341
rect 3130 328 3590 331
rect 2602 318 2990 321
rect 854 303 857 307
rect 853 302 858 303
rect 863 302 864 307
rect 1886 303 1889 307
rect 1885 302 1890 303
rect 1895 302 1896 307
rect 2910 303 2913 307
rect 2909 302 2914 303
rect 2919 302 2920 307
rect 1562 298 1853 301
rect 1902 298 2222 301
rect 2234 298 2438 301
rect 1162 288 1518 291
rect 1902 291 1905 298
rect 1778 288 1905 291
rect 1914 288 2478 291
rect 2530 288 3022 291
rect 482 278 1262 281
rect 1506 278 1934 281
rect 2066 278 2206 281
rect 2458 278 3182 281
rect 298 268 1022 271
rect 1530 268 1582 271
rect 1706 268 1910 271
rect 2474 268 2590 271
rect 3010 268 3174 271
rect 1538 258 1950 261
rect 1970 258 2190 261
rect 3006 261 3009 268
rect 2402 258 3009 261
rect 1538 248 3622 251
rect 1194 238 1838 241
rect 1858 238 2518 241
rect 1442 228 2510 231
rect 1354 218 1622 221
rect 350 203 353 207
rect 349 202 354 203
rect 359 202 360 207
rect 1366 203 1369 207
rect 1365 202 1370 203
rect 1375 202 1376 207
rect 2390 203 2393 207
rect 2389 202 2394 203
rect 2399 202 2400 207
rect 3414 203 3417 207
rect 3413 202 3418 203
rect 3423 202 3424 207
rect 1146 188 2470 191
rect 3006 182 3009 187
rect 1074 178 1590 181
rect 2202 178 2918 181
rect 1658 168 1950 171
rect 2194 168 2702 171
rect 3562 168 3565 171
rect 3578 168 3677 171
rect 3722 168 3741 171
rect 1202 158 1286 161
rect 1402 158 3294 161
rect 3554 158 3558 161
rect 2730 148 2974 151
rect 3162 148 3165 151
rect 3370 148 3678 151
rect 3718 151 3721 158
rect 3718 148 3725 151
rect 2698 138 2838 141
rect 3042 138 3414 141
rect 3706 128 3709 131
rect 854 103 857 107
rect 853 102 858 103
rect 863 102 864 107
rect 1886 103 1889 107
rect 1885 102 1890 103
rect 1895 102 1896 107
rect 2910 103 2913 107
rect 2909 102 2914 103
rect 2919 102 2920 107
rect 3146 78 3181 81
rect 3682 78 3718 81
rect 3758 72 3761 78
rect 514 68 1662 71
rect 3362 68 3469 71
rect 3594 68 3693 71
rect 3482 58 3485 61
rect 3390 42 3393 47
rect 3330 38 3334 41
rect 350 3 353 7
rect 349 2 354 3
rect 359 2 360 7
rect 1366 3 1369 7
rect 1365 2 1370 3
rect 1375 2 1376 7
rect 2390 3 2393 7
rect 2389 2 2394 3
rect 2399 2 2400 7
rect 3414 3 3417 7
rect 3413 2 3418 3
rect 3423 2 3424 7
<< m6contact >>
rect 344 3603 346 3607
rect 346 3603 349 3607
rect 354 3603 357 3607
rect 357 3603 359 3607
rect 344 3602 349 3603
rect 354 3602 359 3603
rect 1360 3603 1362 3607
rect 1362 3603 1365 3607
rect 1370 3603 1373 3607
rect 1373 3603 1375 3607
rect 1360 3602 1365 3603
rect 1370 3602 1375 3603
rect 2384 3603 2386 3607
rect 2386 3603 2389 3607
rect 2394 3603 2397 3607
rect 2397 3603 2399 3607
rect 2384 3602 2389 3603
rect 2394 3602 2399 3603
rect 3408 3603 3410 3607
rect 3410 3603 3413 3607
rect 3418 3603 3421 3607
rect 3421 3603 3423 3607
rect 3408 3602 3413 3603
rect 3418 3602 3423 3603
rect 3565 3547 3570 3552
rect 3613 3537 3618 3542
rect 1805 3527 1810 3532
rect 3741 3527 3746 3532
rect 3501 3517 3506 3522
rect 848 3503 850 3507
rect 850 3503 853 3507
rect 858 3503 861 3507
rect 861 3503 863 3507
rect 848 3502 853 3503
rect 858 3502 863 3503
rect 1880 3503 1882 3507
rect 1882 3503 1885 3507
rect 1890 3503 1893 3507
rect 1893 3503 1895 3507
rect 1880 3502 1885 3503
rect 1890 3502 1895 3503
rect 2904 3503 2906 3507
rect 2906 3503 2909 3507
rect 2914 3503 2917 3507
rect 2917 3503 2919 3507
rect 2904 3502 2909 3503
rect 2914 3502 2919 3503
rect 3741 3457 3746 3462
rect 3597 3437 3602 3442
rect 3661 3437 3666 3442
rect 344 3403 346 3407
rect 346 3403 349 3407
rect 354 3403 357 3407
rect 357 3403 359 3407
rect 344 3402 349 3403
rect 354 3402 359 3403
rect 1360 3403 1362 3407
rect 1362 3403 1365 3407
rect 1370 3403 1373 3407
rect 1373 3403 1375 3407
rect 1360 3402 1365 3403
rect 1370 3402 1375 3403
rect 2384 3403 2386 3407
rect 2386 3403 2389 3407
rect 2394 3403 2397 3407
rect 2397 3403 2399 3407
rect 2384 3402 2389 3403
rect 2394 3402 2399 3403
rect 3408 3403 3410 3407
rect 3410 3403 3413 3407
rect 3418 3403 3421 3407
rect 3421 3403 3423 3407
rect 3408 3402 3413 3403
rect 3418 3402 3423 3403
rect 848 3303 850 3307
rect 850 3303 853 3307
rect 858 3303 861 3307
rect 861 3303 863 3307
rect 848 3302 853 3303
rect 858 3302 863 3303
rect 1880 3303 1882 3307
rect 1882 3303 1885 3307
rect 1890 3303 1893 3307
rect 1893 3303 1895 3307
rect 1880 3302 1885 3303
rect 1890 3302 1895 3303
rect 2904 3303 2906 3307
rect 2906 3303 2909 3307
rect 2914 3303 2917 3307
rect 2917 3303 2919 3307
rect 2904 3302 2909 3303
rect 2914 3302 2919 3303
rect 344 3203 346 3207
rect 346 3203 349 3207
rect 354 3203 357 3207
rect 357 3203 359 3207
rect 344 3202 349 3203
rect 354 3202 359 3203
rect 1360 3203 1362 3207
rect 1362 3203 1365 3207
rect 1370 3203 1373 3207
rect 1373 3203 1375 3207
rect 1360 3202 1365 3203
rect 1370 3202 1375 3203
rect 2384 3203 2386 3207
rect 2386 3203 2389 3207
rect 2394 3203 2397 3207
rect 2397 3203 2399 3207
rect 2384 3202 2389 3203
rect 2394 3202 2399 3203
rect 3408 3203 3410 3207
rect 3410 3203 3413 3207
rect 3418 3203 3421 3207
rect 3421 3203 3423 3207
rect 3408 3202 3413 3203
rect 3418 3202 3423 3203
rect 848 3103 850 3107
rect 850 3103 853 3107
rect 858 3103 861 3107
rect 861 3103 863 3107
rect 848 3102 853 3103
rect 858 3102 863 3103
rect 1880 3103 1882 3107
rect 1882 3103 1885 3107
rect 1890 3103 1893 3107
rect 1893 3103 1895 3107
rect 1880 3102 1885 3103
rect 1890 3102 1895 3103
rect 2904 3103 2906 3107
rect 2906 3103 2909 3107
rect 2914 3103 2917 3107
rect 2917 3103 2919 3107
rect 2904 3102 2909 3103
rect 2914 3102 2919 3103
rect 3581 3087 3586 3092
rect 3645 3087 3650 3092
rect 3709 3087 3714 3092
rect 3693 3077 3698 3082
rect 3725 3077 3730 3082
rect 344 3003 346 3007
rect 346 3003 349 3007
rect 354 3003 357 3007
rect 357 3003 359 3007
rect 344 3002 349 3003
rect 354 3002 359 3003
rect 1360 3003 1362 3007
rect 1362 3003 1365 3007
rect 1370 3003 1373 3007
rect 1373 3003 1375 3007
rect 1360 3002 1365 3003
rect 1370 3002 1375 3003
rect 2384 3003 2386 3007
rect 2386 3003 2389 3007
rect 2394 3003 2397 3007
rect 2397 3003 2399 3007
rect 2384 3002 2389 3003
rect 2394 3002 2399 3003
rect 3408 3003 3410 3007
rect 3410 3003 3413 3007
rect 3418 3003 3421 3007
rect 3421 3003 3423 3007
rect 3408 3002 3413 3003
rect 3418 3002 3423 3003
rect 848 2903 850 2907
rect 850 2903 853 2907
rect 858 2903 861 2907
rect 861 2903 863 2907
rect 848 2902 853 2903
rect 858 2902 863 2903
rect 1880 2903 1882 2907
rect 1882 2903 1885 2907
rect 1890 2903 1893 2907
rect 1893 2903 1895 2907
rect 1880 2902 1885 2903
rect 1890 2902 1895 2903
rect 2904 2903 2906 2907
rect 2906 2903 2909 2907
rect 2914 2903 2917 2907
rect 2917 2903 2919 2907
rect 2904 2902 2909 2903
rect 2914 2902 2919 2903
rect 344 2803 346 2807
rect 346 2803 349 2807
rect 354 2803 357 2807
rect 357 2803 359 2807
rect 344 2802 349 2803
rect 354 2802 359 2803
rect 1360 2803 1362 2807
rect 1362 2803 1365 2807
rect 1370 2803 1373 2807
rect 1373 2803 1375 2807
rect 1360 2802 1365 2803
rect 1370 2802 1375 2803
rect 2384 2803 2386 2807
rect 2386 2803 2389 2807
rect 2394 2803 2397 2807
rect 2397 2803 2399 2807
rect 2384 2802 2389 2803
rect 2394 2802 2399 2803
rect 3408 2803 3410 2807
rect 3410 2803 3413 2807
rect 3418 2803 3421 2807
rect 3421 2803 3423 2807
rect 3408 2802 3413 2803
rect 3418 2802 3423 2803
rect 1789 2797 1794 2802
rect 3453 2747 3458 2752
rect 1805 2727 1810 2732
rect 848 2703 850 2707
rect 850 2703 853 2707
rect 858 2703 861 2707
rect 861 2703 863 2707
rect 848 2702 853 2703
rect 858 2702 863 2703
rect 1880 2703 1882 2707
rect 1882 2703 1885 2707
rect 1890 2703 1893 2707
rect 1893 2703 1895 2707
rect 1880 2702 1885 2703
rect 1890 2702 1895 2703
rect 2904 2703 2906 2707
rect 2906 2703 2909 2707
rect 2914 2703 2917 2707
rect 2917 2703 2919 2707
rect 2904 2702 2909 2703
rect 2914 2702 2919 2703
rect 344 2603 346 2607
rect 346 2603 349 2607
rect 354 2603 357 2607
rect 357 2603 359 2607
rect 344 2602 349 2603
rect 354 2602 359 2603
rect 1360 2603 1362 2607
rect 1362 2603 1365 2607
rect 1370 2603 1373 2607
rect 1373 2603 1375 2607
rect 1360 2602 1365 2603
rect 1370 2602 1375 2603
rect 2384 2603 2386 2607
rect 2386 2603 2389 2607
rect 2394 2603 2397 2607
rect 2397 2603 2399 2607
rect 2384 2602 2389 2603
rect 2394 2602 2399 2603
rect 3408 2603 3410 2607
rect 3410 2603 3413 2607
rect 3418 2603 3421 2607
rect 3421 2603 3423 2607
rect 3408 2602 3413 2603
rect 3418 2602 3423 2603
rect 3181 2537 3186 2542
rect 3725 2537 3730 2542
rect 848 2503 850 2507
rect 850 2503 853 2507
rect 858 2503 861 2507
rect 861 2503 863 2507
rect 848 2502 853 2503
rect 858 2502 863 2503
rect 1880 2503 1882 2507
rect 1882 2503 1885 2507
rect 1890 2503 1893 2507
rect 1893 2503 1895 2507
rect 1880 2502 1885 2503
rect 1890 2502 1895 2503
rect 2904 2503 2906 2507
rect 2906 2503 2909 2507
rect 2914 2503 2917 2507
rect 2917 2503 2919 2507
rect 2904 2502 2909 2503
rect 2914 2502 2919 2503
rect 3469 2417 3474 2422
rect 344 2403 346 2407
rect 346 2403 349 2407
rect 354 2403 357 2407
rect 357 2403 359 2407
rect 344 2402 349 2403
rect 354 2402 359 2403
rect 1360 2403 1362 2407
rect 1362 2403 1365 2407
rect 1370 2403 1373 2407
rect 1373 2403 1375 2407
rect 1360 2402 1365 2403
rect 1370 2402 1375 2403
rect 2384 2403 2386 2407
rect 2386 2403 2389 2407
rect 2394 2403 2397 2407
rect 2397 2403 2399 2407
rect 2384 2402 2389 2403
rect 2394 2402 2399 2403
rect 3408 2403 3410 2407
rect 3410 2403 3413 2407
rect 3418 2403 3421 2407
rect 3421 2403 3423 2407
rect 3408 2402 3413 2403
rect 3418 2402 3423 2403
rect 3629 2367 3634 2372
rect 848 2303 850 2307
rect 850 2303 853 2307
rect 858 2303 861 2307
rect 861 2303 863 2307
rect 848 2302 853 2303
rect 858 2302 863 2303
rect 1880 2303 1882 2307
rect 1882 2303 1885 2307
rect 1890 2303 1893 2307
rect 1893 2303 1895 2307
rect 1880 2302 1885 2303
rect 1890 2302 1895 2303
rect 2904 2303 2906 2307
rect 2906 2303 2909 2307
rect 2914 2303 2917 2307
rect 2917 2303 2919 2307
rect 2904 2302 2909 2303
rect 2914 2302 2919 2303
rect 2893 2297 2898 2302
rect 3677 2287 3682 2292
rect 1485 2277 1490 2282
rect 1509 2267 1514 2272
rect 2893 2267 2898 2272
rect 3693 2277 3698 2282
rect 3517 2247 3522 2252
rect 344 2203 346 2207
rect 346 2203 349 2207
rect 354 2203 357 2207
rect 357 2203 359 2207
rect 344 2202 349 2203
rect 354 2202 359 2203
rect 1360 2203 1362 2207
rect 1362 2203 1365 2207
rect 1370 2203 1373 2207
rect 1373 2203 1375 2207
rect 1360 2202 1365 2203
rect 1370 2202 1375 2203
rect 2384 2203 2386 2207
rect 2386 2203 2389 2207
rect 2394 2203 2397 2207
rect 2397 2203 2399 2207
rect 2384 2202 2389 2203
rect 2394 2202 2399 2203
rect 3408 2203 3410 2207
rect 3410 2203 3413 2207
rect 3418 2203 3421 2207
rect 3421 2203 3423 2207
rect 3408 2202 3413 2203
rect 3418 2202 3423 2203
rect 3661 2137 3666 2142
rect 848 2103 850 2107
rect 850 2103 853 2107
rect 858 2103 861 2107
rect 861 2103 863 2107
rect 848 2102 853 2103
rect 858 2102 863 2103
rect 1880 2103 1882 2107
rect 1882 2103 1885 2107
rect 1890 2103 1893 2107
rect 1893 2103 1895 2107
rect 1880 2102 1885 2103
rect 1890 2102 1895 2103
rect 2904 2103 2906 2107
rect 2906 2103 2909 2107
rect 2914 2103 2917 2107
rect 2917 2103 2919 2107
rect 2904 2102 2909 2103
rect 2914 2102 2919 2103
rect 3533 2077 3538 2082
rect 3661 2057 3666 2062
rect 1789 2047 1794 2052
rect 3693 2047 3698 2052
rect 3709 2047 3714 2052
rect 3709 2037 3714 2042
rect 3437 2027 3442 2032
rect 344 2003 346 2007
rect 346 2003 349 2007
rect 354 2003 357 2007
rect 357 2003 359 2007
rect 344 2002 349 2003
rect 354 2002 359 2003
rect 1360 2003 1362 2007
rect 1362 2003 1365 2007
rect 1370 2003 1373 2007
rect 1373 2003 1375 2007
rect 1360 2002 1365 2003
rect 1370 2002 1375 2003
rect 2384 2003 2386 2007
rect 2386 2003 2389 2007
rect 2394 2003 2397 2007
rect 2397 2003 2399 2007
rect 2384 2002 2389 2003
rect 2394 2002 2399 2003
rect 3408 2003 3410 2007
rect 3410 2003 3413 2007
rect 3418 2003 3421 2007
rect 3421 2003 3423 2007
rect 3408 2002 3413 2003
rect 3418 2002 3423 2003
rect 3613 1947 3618 1952
rect 3133 1937 3138 1942
rect 3757 1937 3762 1942
rect 3613 1927 3618 1932
rect 848 1903 850 1907
rect 850 1903 853 1907
rect 858 1903 861 1907
rect 861 1903 863 1907
rect 848 1902 853 1903
rect 858 1902 863 1903
rect 1880 1903 1882 1907
rect 1882 1903 1885 1907
rect 1890 1903 1893 1907
rect 1893 1903 1895 1907
rect 1880 1902 1885 1903
rect 1890 1902 1895 1903
rect 2904 1903 2906 1907
rect 2906 1903 2909 1907
rect 2914 1903 2917 1907
rect 2917 1903 2919 1907
rect 2904 1902 2909 1903
rect 2914 1902 2919 1903
rect 3773 1867 3778 1872
rect 3565 1837 3570 1842
rect 2813 1817 2818 1822
rect 344 1803 346 1807
rect 346 1803 349 1807
rect 354 1803 357 1807
rect 357 1803 359 1807
rect 344 1802 349 1803
rect 354 1802 359 1803
rect 1360 1803 1362 1807
rect 1362 1803 1365 1807
rect 1370 1803 1373 1807
rect 1373 1803 1375 1807
rect 1360 1802 1365 1803
rect 1370 1802 1375 1803
rect 2384 1803 2386 1807
rect 2386 1803 2389 1807
rect 2394 1803 2397 1807
rect 2397 1803 2399 1807
rect 2384 1802 2389 1803
rect 2394 1802 2399 1803
rect 3408 1803 3410 1807
rect 3410 1803 3413 1807
rect 3418 1803 3421 1807
rect 3421 1803 3423 1807
rect 3408 1802 3413 1803
rect 3418 1802 3423 1803
rect 3581 1757 3586 1762
rect 3373 1747 3378 1752
rect 3725 1727 3730 1732
rect 848 1703 850 1707
rect 850 1703 853 1707
rect 858 1703 861 1707
rect 861 1703 863 1707
rect 848 1702 853 1703
rect 858 1702 863 1703
rect 1880 1703 1882 1707
rect 1882 1703 1885 1707
rect 1890 1703 1893 1707
rect 1893 1703 1895 1707
rect 1880 1702 1885 1703
rect 1890 1702 1895 1703
rect 2904 1703 2906 1707
rect 2906 1703 2909 1707
rect 2914 1703 2917 1707
rect 2917 1703 2919 1707
rect 2904 1702 2909 1703
rect 2914 1702 2919 1703
rect 3549 1687 3554 1692
rect 3709 1637 3714 1642
rect 3565 1607 3570 1612
rect 344 1603 346 1607
rect 346 1603 349 1607
rect 354 1603 357 1607
rect 357 1603 359 1607
rect 344 1602 349 1603
rect 354 1602 359 1603
rect 1360 1603 1362 1607
rect 1362 1603 1365 1607
rect 1370 1603 1373 1607
rect 1373 1603 1375 1607
rect 1360 1602 1365 1603
rect 1370 1602 1375 1603
rect 2384 1603 2386 1607
rect 2386 1603 2389 1607
rect 2394 1603 2397 1607
rect 2397 1603 2399 1607
rect 2384 1602 2389 1603
rect 2394 1602 2399 1603
rect 3408 1603 3410 1607
rect 3410 1603 3413 1607
rect 3418 1603 3421 1607
rect 3421 1603 3423 1607
rect 3408 1602 3413 1603
rect 3418 1602 3423 1603
rect 3741 1597 3746 1602
rect 3133 1567 3138 1572
rect 1581 1547 1586 1552
rect 3709 1557 3714 1562
rect 3533 1547 3538 1552
rect 3501 1537 3506 1542
rect 3533 1537 3538 1542
rect 3677 1507 3682 1512
rect 848 1503 850 1507
rect 850 1503 853 1507
rect 858 1503 861 1507
rect 861 1503 863 1507
rect 848 1502 853 1503
rect 858 1502 863 1503
rect 1880 1503 1882 1507
rect 1882 1503 1885 1507
rect 1890 1503 1893 1507
rect 1893 1503 1895 1507
rect 1880 1502 1885 1503
rect 1890 1502 1895 1503
rect 2904 1503 2906 1507
rect 2906 1503 2909 1507
rect 2914 1503 2917 1507
rect 2917 1503 2919 1507
rect 2904 1502 2909 1503
rect 2914 1502 2919 1503
rect 3485 1487 3490 1492
rect 3677 1487 3682 1492
rect 3693 1477 3698 1482
rect 3629 1457 3634 1462
rect 3597 1447 3602 1452
rect 3629 1447 3634 1452
rect 344 1403 346 1407
rect 346 1403 349 1407
rect 354 1403 357 1407
rect 357 1403 359 1407
rect 344 1402 349 1403
rect 354 1402 359 1403
rect 1360 1403 1362 1407
rect 1362 1403 1365 1407
rect 1370 1403 1373 1407
rect 1373 1403 1375 1407
rect 1360 1402 1365 1403
rect 1370 1402 1375 1403
rect 2384 1403 2386 1407
rect 2386 1403 2389 1407
rect 2394 1403 2397 1407
rect 2397 1403 2399 1407
rect 2384 1402 2389 1403
rect 2394 1402 2399 1403
rect 3408 1403 3410 1407
rect 3410 1403 3413 1407
rect 3418 1403 3421 1407
rect 3421 1403 3423 1407
rect 3408 1402 3413 1403
rect 3418 1402 3423 1403
rect 3325 1387 3330 1392
rect 3597 1377 3602 1382
rect 3645 1377 3650 1382
rect 3693 1367 3698 1372
rect 3645 1357 3650 1362
rect 3501 1327 3506 1332
rect 3725 1327 3730 1332
rect 3629 1317 3634 1322
rect 3149 1307 3154 1312
rect 848 1303 850 1307
rect 850 1303 853 1307
rect 858 1303 861 1307
rect 861 1303 863 1307
rect 848 1302 853 1303
rect 858 1302 863 1303
rect 1880 1303 1882 1307
rect 1882 1303 1885 1307
rect 1890 1303 1893 1307
rect 1893 1303 1895 1307
rect 1880 1302 1885 1303
rect 1890 1302 1895 1303
rect 2904 1303 2906 1307
rect 2906 1303 2909 1307
rect 2914 1303 2917 1307
rect 2917 1303 2919 1307
rect 2904 1302 2909 1303
rect 2914 1302 2919 1303
rect 3069 1277 3074 1282
rect 3645 1277 3650 1282
rect 3533 1267 3538 1272
rect 3645 1257 3650 1262
rect 3757 1247 3762 1252
rect 3005 1217 3010 1222
rect 344 1203 346 1207
rect 346 1203 349 1207
rect 354 1203 357 1207
rect 357 1203 359 1207
rect 344 1202 349 1203
rect 354 1202 359 1203
rect 1360 1203 1362 1207
rect 1362 1203 1365 1207
rect 1370 1203 1373 1207
rect 1373 1203 1375 1207
rect 1360 1202 1365 1203
rect 1370 1202 1375 1203
rect 2384 1203 2386 1207
rect 2386 1203 2389 1207
rect 2394 1203 2397 1207
rect 2397 1203 2399 1207
rect 2384 1202 2389 1203
rect 2394 1202 2399 1203
rect 3408 1203 3410 1207
rect 3410 1203 3413 1207
rect 3418 1203 3421 1207
rect 3421 1203 3423 1207
rect 3408 1202 3413 1203
rect 3418 1202 3423 1203
rect 3757 1197 3762 1202
rect 3453 1157 3458 1162
rect 3533 1147 3538 1152
rect 3389 1137 3394 1142
rect 3581 1117 3586 1122
rect 848 1103 850 1107
rect 850 1103 853 1107
rect 858 1103 861 1107
rect 861 1103 863 1107
rect 848 1102 853 1103
rect 858 1102 863 1103
rect 1880 1103 1882 1107
rect 1882 1103 1885 1107
rect 1890 1103 1893 1107
rect 1893 1103 1895 1107
rect 1880 1102 1885 1103
rect 1890 1102 1895 1103
rect 2904 1103 2906 1107
rect 2906 1103 2909 1107
rect 2914 1103 2917 1107
rect 2917 1103 2919 1107
rect 2904 1102 2909 1103
rect 2914 1102 2919 1103
rect 3037 1097 3042 1102
rect 1597 1067 1602 1072
rect 3773 1067 3778 1072
rect 3373 1047 3378 1052
rect 3029 1007 3034 1012
rect 344 1003 346 1007
rect 346 1003 349 1007
rect 354 1003 357 1007
rect 357 1003 359 1007
rect 344 1002 349 1003
rect 354 1002 359 1003
rect 1360 1003 1362 1007
rect 1362 1003 1365 1007
rect 1370 1003 1373 1007
rect 1373 1003 1375 1007
rect 1360 1002 1365 1003
rect 1370 1002 1375 1003
rect 2384 1003 2386 1007
rect 2386 1003 2389 1007
rect 2394 1003 2397 1007
rect 2397 1003 2399 1007
rect 2384 1002 2389 1003
rect 2394 1002 2399 1003
rect 3408 1003 3410 1007
rect 3410 1003 3413 1007
rect 3418 1003 3421 1007
rect 3421 1003 3423 1007
rect 3408 1002 3413 1003
rect 3418 1002 3423 1003
rect 3613 997 3618 1002
rect 3613 987 3618 992
rect 2877 947 2882 952
rect 2877 927 2882 932
rect 3629 917 3634 922
rect 848 903 850 907
rect 850 903 853 907
rect 858 903 861 907
rect 861 903 863 907
rect 848 902 853 903
rect 858 902 863 903
rect 1880 903 1882 907
rect 1882 903 1885 907
rect 1890 903 1893 907
rect 1893 903 1895 907
rect 1880 902 1885 903
rect 1890 902 1895 903
rect 2904 903 2906 907
rect 2906 903 2909 907
rect 2914 903 2917 907
rect 2917 903 2919 907
rect 2904 902 2909 903
rect 2914 902 2919 903
rect 344 803 346 807
rect 346 803 349 807
rect 354 803 357 807
rect 357 803 359 807
rect 344 802 349 803
rect 354 802 359 803
rect 1360 803 1362 807
rect 1362 803 1365 807
rect 1370 803 1373 807
rect 1373 803 1375 807
rect 1360 802 1365 803
rect 1370 802 1375 803
rect 2384 803 2386 807
rect 2386 803 2389 807
rect 2394 803 2397 807
rect 2397 803 2399 807
rect 2384 802 2389 803
rect 2394 802 2399 803
rect 3408 803 3410 807
rect 3410 803 3413 807
rect 3418 803 3421 807
rect 3421 803 3423 807
rect 3408 802 3413 803
rect 3418 802 3423 803
rect 3725 777 3730 782
rect 3437 747 3442 752
rect 3613 737 3618 742
rect 848 703 850 707
rect 850 703 853 707
rect 858 703 861 707
rect 861 703 863 707
rect 848 702 853 703
rect 858 702 863 703
rect 1880 703 1882 707
rect 1882 703 1885 707
rect 1890 703 1893 707
rect 1893 703 1895 707
rect 1880 702 1885 703
rect 1890 702 1895 703
rect 2904 703 2906 707
rect 2906 703 2909 707
rect 2914 703 2917 707
rect 2917 703 2919 707
rect 2904 702 2909 703
rect 2914 702 2919 703
rect 3165 697 3170 702
rect 3533 687 3538 692
rect 1597 667 1602 672
rect 3149 657 3154 662
rect 3645 637 3650 642
rect 344 603 346 607
rect 346 603 349 607
rect 354 603 357 607
rect 357 603 359 607
rect 344 602 349 603
rect 354 602 359 603
rect 1360 603 1362 607
rect 1362 603 1365 607
rect 1370 603 1373 607
rect 1373 603 1375 607
rect 1360 602 1365 603
rect 1370 602 1375 603
rect 2384 603 2386 607
rect 2386 603 2389 607
rect 2394 603 2397 607
rect 2397 603 2399 607
rect 2384 602 2389 603
rect 2394 602 2399 603
rect 3408 603 3410 607
rect 3410 603 3413 607
rect 3418 603 3421 607
rect 3421 603 3423 607
rect 3408 602 3413 603
rect 3418 602 3423 603
rect 2749 577 2754 582
rect 1581 547 1586 552
rect 3069 507 3074 512
rect 848 503 850 507
rect 850 503 853 507
rect 858 503 861 507
rect 861 503 863 507
rect 848 502 853 503
rect 858 502 863 503
rect 1880 503 1882 507
rect 1882 503 1885 507
rect 1890 503 1893 507
rect 1893 503 1895 507
rect 1880 502 1885 503
rect 1890 502 1895 503
rect 2904 503 2906 507
rect 2906 503 2909 507
rect 2914 503 2917 507
rect 2917 503 2919 507
rect 2904 502 2909 503
rect 2914 502 2919 503
rect 2813 457 2818 462
rect 2749 447 2754 452
rect 3517 427 3522 432
rect 344 403 346 407
rect 346 403 349 407
rect 354 403 357 407
rect 357 403 359 407
rect 344 402 349 403
rect 354 402 359 403
rect 1360 403 1362 407
rect 1362 403 1365 407
rect 1370 403 1373 407
rect 1373 403 1375 407
rect 1360 402 1365 403
rect 1370 402 1375 403
rect 2384 403 2386 407
rect 2386 403 2389 407
rect 2394 403 2397 407
rect 2397 403 2399 407
rect 2384 402 2389 403
rect 2394 402 2399 403
rect 3408 403 3410 407
rect 3410 403 3413 407
rect 3418 403 3421 407
rect 3421 403 3423 407
rect 3408 402 3413 403
rect 3418 402 3423 403
rect 3629 367 3634 372
rect 3661 357 3666 362
rect 3501 347 3506 352
rect 3597 347 3602 352
rect 3581 337 3586 342
rect 848 303 850 307
rect 850 303 853 307
rect 858 303 861 307
rect 861 303 863 307
rect 848 302 853 303
rect 858 302 863 303
rect 1880 303 1882 307
rect 1882 303 1885 307
rect 1890 303 1893 307
rect 1893 303 1895 307
rect 1880 302 1885 303
rect 1890 302 1895 303
rect 2904 303 2906 307
rect 2906 303 2909 307
rect 2914 303 2917 307
rect 2917 303 2919 307
rect 2904 302 2909 303
rect 2914 302 2919 303
rect 1853 297 1858 302
rect 1853 237 1858 242
rect 344 203 346 207
rect 346 203 349 207
rect 354 203 357 207
rect 357 203 359 207
rect 344 202 349 203
rect 354 202 359 203
rect 1360 203 1362 207
rect 1362 203 1365 207
rect 1370 203 1373 207
rect 1373 203 1375 207
rect 1360 202 1365 203
rect 1370 202 1375 203
rect 2384 203 2386 207
rect 2386 203 2389 207
rect 2394 203 2397 207
rect 2397 203 2399 207
rect 2384 202 2389 203
rect 2394 202 2399 203
rect 3408 203 3410 207
rect 3410 203 3413 207
rect 3418 203 3421 207
rect 3421 203 3423 207
rect 3408 202 3413 203
rect 3418 202 3423 203
rect 3005 187 3010 192
rect 3565 167 3570 172
rect 3677 167 3682 172
rect 3741 167 3746 172
rect 3549 157 3554 162
rect 3165 147 3170 152
rect 3725 147 3730 152
rect 3709 127 3714 132
rect 848 103 850 107
rect 850 103 853 107
rect 858 103 861 107
rect 861 103 863 107
rect 848 102 853 103
rect 858 102 863 103
rect 1880 103 1882 107
rect 1882 103 1885 107
rect 1890 103 1893 107
rect 1893 103 1895 107
rect 1880 102 1885 103
rect 1890 102 1895 103
rect 2904 103 2906 107
rect 2906 103 2909 107
rect 2914 103 2917 107
rect 2917 103 2919 107
rect 2904 102 2909 103
rect 2914 102 2919 103
rect 3181 77 3186 82
rect 3677 77 3682 82
rect 3469 67 3474 72
rect 3693 67 3698 72
rect 3757 67 3762 72
rect 3485 57 3490 62
rect 3389 47 3394 52
rect 3325 37 3330 42
rect 344 3 346 7
rect 346 3 349 7
rect 354 3 357 7
rect 357 3 359 7
rect 344 2 349 3
rect 354 2 359 3
rect 1360 3 1362 7
rect 1362 3 1365 7
rect 1370 3 1373 7
rect 1373 3 1375 7
rect 1360 2 1365 3
rect 1370 2 1375 3
rect 2384 3 2386 7
rect 2386 3 2389 7
rect 2394 3 2397 7
rect 2397 3 2399 7
rect 2384 2 2389 3
rect 2394 2 2399 3
rect 3408 3 3410 7
rect 3410 3 3413 7
rect 3418 3 3421 7
rect 3421 3 3423 7
rect 3408 2 3413 3
rect 3418 2 3423 3
<< metal6 >>
rect 344 3607 360 3630
rect 349 3602 354 3607
rect 359 3602 360 3607
rect 344 3407 360 3602
rect 349 3402 354 3407
rect 359 3402 360 3407
rect 344 3207 360 3402
rect 349 3202 354 3207
rect 359 3202 360 3207
rect 344 3007 360 3202
rect 349 3002 354 3007
rect 359 3002 360 3007
rect 344 2807 360 3002
rect 349 2802 354 2807
rect 359 2802 360 2807
rect 344 2607 360 2802
rect 349 2602 354 2607
rect 359 2602 360 2607
rect 344 2407 360 2602
rect 349 2402 354 2407
rect 359 2402 360 2407
rect 344 2207 360 2402
rect 349 2202 354 2207
rect 359 2202 360 2207
rect 344 2007 360 2202
rect 349 2002 354 2007
rect 359 2002 360 2007
rect 344 1807 360 2002
rect 349 1802 354 1807
rect 359 1802 360 1807
rect 344 1607 360 1802
rect 349 1602 354 1607
rect 359 1602 360 1607
rect 344 1407 360 1602
rect 349 1402 354 1407
rect 359 1402 360 1407
rect 344 1207 360 1402
rect 349 1202 354 1207
rect 359 1202 360 1207
rect 344 1007 360 1202
rect 349 1002 354 1007
rect 359 1002 360 1007
rect 344 807 360 1002
rect 349 802 354 807
rect 359 802 360 807
rect 344 607 360 802
rect 349 602 354 607
rect 359 602 360 607
rect 344 407 360 602
rect 349 402 354 407
rect 359 402 360 407
rect 344 207 360 402
rect 349 202 354 207
rect 359 202 360 207
rect 344 7 360 202
rect 349 2 354 7
rect 359 2 360 7
rect 344 -30 360 2
rect 848 3507 864 3630
rect 853 3502 858 3507
rect 863 3502 864 3507
rect 848 3307 864 3502
rect 853 3302 858 3307
rect 863 3302 864 3307
rect 848 3107 864 3302
rect 853 3102 858 3107
rect 863 3102 864 3107
rect 848 2907 864 3102
rect 853 2902 858 2907
rect 863 2902 864 2907
rect 848 2707 864 2902
rect 853 2702 858 2707
rect 863 2702 864 2707
rect 848 2507 864 2702
rect 853 2502 858 2507
rect 863 2502 864 2507
rect 848 2307 864 2502
rect 853 2302 858 2307
rect 863 2302 864 2307
rect 848 2107 864 2302
rect 853 2102 858 2107
rect 863 2102 864 2107
rect 848 1907 864 2102
rect 853 1902 858 1907
rect 863 1902 864 1907
rect 848 1707 864 1902
rect 853 1702 858 1707
rect 863 1702 864 1707
rect 848 1507 864 1702
rect 853 1502 858 1507
rect 863 1502 864 1507
rect 848 1307 864 1502
rect 853 1302 858 1307
rect 863 1302 864 1307
rect 848 1107 864 1302
rect 853 1102 858 1107
rect 863 1102 864 1107
rect 848 907 864 1102
rect 853 902 858 907
rect 863 902 864 907
rect 848 707 864 902
rect 853 702 858 707
rect 863 702 864 707
rect 848 507 864 702
rect 853 502 858 507
rect 863 502 864 507
rect 848 307 864 502
rect 853 302 858 307
rect 863 302 864 307
rect 848 107 864 302
rect 853 102 858 107
rect 863 102 864 107
rect 848 -30 864 102
rect 1360 3607 1376 3630
rect 1365 3602 1370 3607
rect 1375 3602 1376 3607
rect 1360 3407 1376 3602
rect 1365 3402 1370 3407
rect 1375 3402 1376 3407
rect 1360 3207 1376 3402
rect 1365 3202 1370 3207
rect 1375 3202 1376 3207
rect 1360 3007 1376 3202
rect 1365 3002 1370 3007
rect 1375 3002 1376 3007
rect 1360 2807 1376 3002
rect 1365 2802 1370 2807
rect 1375 2802 1376 2807
rect 1360 2607 1376 2802
rect 1365 2602 1370 2607
rect 1375 2602 1376 2607
rect 1360 2407 1376 2602
rect 1365 2402 1370 2407
rect 1375 2402 1376 2407
rect 1360 2207 1376 2402
rect 1485 2272 1490 2277
rect 1485 2267 1509 2272
rect 1365 2202 1370 2207
rect 1375 2202 1376 2207
rect 1360 2007 1376 2202
rect 1789 2052 1794 2797
rect 1805 2732 1810 3527
rect 1880 3507 1896 3630
rect 1885 3502 1890 3507
rect 1895 3502 1896 3507
rect 1880 3307 1896 3502
rect 1885 3302 1890 3307
rect 1895 3302 1896 3307
rect 1880 3107 1896 3302
rect 1885 3102 1890 3107
rect 1895 3102 1896 3107
rect 1880 2907 1896 3102
rect 1885 2902 1890 2907
rect 1895 2902 1896 2907
rect 1880 2707 1896 2902
rect 1885 2702 1890 2707
rect 1895 2702 1896 2707
rect 1880 2507 1896 2702
rect 1885 2502 1890 2507
rect 1895 2502 1896 2507
rect 1880 2307 1896 2502
rect 1885 2302 1890 2307
rect 1895 2302 1896 2307
rect 1880 2107 1896 2302
rect 1885 2102 1890 2107
rect 1895 2102 1896 2107
rect 1365 2002 1370 2007
rect 1375 2002 1376 2007
rect 1360 1807 1376 2002
rect 1365 1802 1370 1807
rect 1375 1802 1376 1807
rect 1360 1607 1376 1802
rect 1365 1602 1370 1607
rect 1375 1602 1376 1607
rect 1360 1407 1376 1602
rect 1880 1907 1896 2102
rect 1885 1902 1890 1907
rect 1895 1902 1896 1907
rect 1880 1707 1896 1902
rect 1885 1702 1890 1707
rect 1895 1702 1896 1707
rect 1365 1402 1370 1407
rect 1375 1402 1376 1407
rect 1360 1207 1376 1402
rect 1365 1202 1370 1207
rect 1375 1202 1376 1207
rect 1360 1007 1376 1202
rect 1365 1002 1370 1007
rect 1375 1002 1376 1007
rect 1360 807 1376 1002
rect 1365 802 1370 807
rect 1375 802 1376 807
rect 1360 607 1376 802
rect 1365 602 1370 607
rect 1375 602 1376 607
rect 1360 407 1376 602
rect 1581 552 1586 1547
rect 1880 1507 1896 1702
rect 1885 1502 1890 1507
rect 1895 1502 1896 1507
rect 1880 1307 1896 1502
rect 1885 1302 1890 1307
rect 1895 1302 1896 1307
rect 1880 1107 1896 1302
rect 1885 1102 1890 1107
rect 1895 1102 1896 1107
rect 1597 672 1602 1067
rect 1880 907 1896 1102
rect 1885 902 1890 907
rect 1895 902 1896 907
rect 1880 707 1896 902
rect 1885 702 1890 707
rect 1895 702 1896 707
rect 1365 402 1370 407
rect 1375 402 1376 407
rect 1360 207 1376 402
rect 1880 507 1896 702
rect 1885 502 1890 507
rect 1895 502 1896 507
rect 1880 307 1896 502
rect 1885 302 1890 307
rect 1895 302 1896 307
rect 1853 242 1858 297
rect 1365 202 1370 207
rect 1375 202 1376 207
rect 1360 7 1376 202
rect 1365 2 1370 7
rect 1375 2 1376 7
rect 1360 -30 1376 2
rect 1880 107 1896 302
rect 1885 102 1890 107
rect 1895 102 1896 107
rect 1880 -30 1896 102
rect 2384 3607 2400 3630
rect 2389 3602 2394 3607
rect 2399 3602 2400 3607
rect 2384 3407 2400 3602
rect 2389 3402 2394 3407
rect 2399 3402 2400 3407
rect 2384 3207 2400 3402
rect 2389 3202 2394 3207
rect 2399 3202 2400 3207
rect 2384 3007 2400 3202
rect 2389 3002 2394 3007
rect 2399 3002 2400 3007
rect 2384 2807 2400 3002
rect 2389 2802 2394 2807
rect 2399 2802 2400 2807
rect 2384 2607 2400 2802
rect 2389 2602 2394 2607
rect 2399 2602 2400 2607
rect 2384 2407 2400 2602
rect 2389 2402 2394 2407
rect 2399 2402 2400 2407
rect 2384 2207 2400 2402
rect 2904 3507 2920 3630
rect 2909 3502 2914 3507
rect 2919 3502 2920 3507
rect 2904 3307 2920 3502
rect 2909 3302 2914 3307
rect 2919 3302 2920 3307
rect 2904 3107 2920 3302
rect 2909 3102 2914 3107
rect 2919 3102 2920 3107
rect 2904 2907 2920 3102
rect 2909 2902 2914 2907
rect 2919 2902 2920 2907
rect 2904 2707 2920 2902
rect 2909 2702 2914 2707
rect 2919 2702 2920 2707
rect 2904 2507 2920 2702
rect 3408 3607 3424 3630
rect 3413 3602 3418 3607
rect 3423 3602 3424 3607
rect 3408 3407 3424 3602
rect 3413 3402 3418 3407
rect 3423 3402 3424 3407
rect 3408 3207 3424 3402
rect 3413 3202 3418 3207
rect 3423 3202 3424 3207
rect 3408 3007 3424 3202
rect 3413 3002 3418 3007
rect 3423 3002 3424 3007
rect 3408 2807 3424 3002
rect 3413 2802 3418 2807
rect 3423 2802 3424 2807
rect 3408 2607 3424 2802
rect 3413 2602 3418 2607
rect 3423 2602 3424 2607
rect 2909 2502 2914 2507
rect 2919 2502 2920 2507
rect 2904 2307 2920 2502
rect 2909 2302 2914 2307
rect 2919 2302 2920 2307
rect 2893 2272 2898 2297
rect 2389 2202 2394 2207
rect 2399 2202 2400 2207
rect 2384 2007 2400 2202
rect 2389 2002 2394 2007
rect 2399 2002 2400 2007
rect 2384 1807 2400 2002
rect 2904 2107 2920 2302
rect 2909 2102 2914 2107
rect 2919 2102 2920 2107
rect 2904 1907 2920 2102
rect 2909 1902 2914 1907
rect 2919 1902 2920 1907
rect 2389 1802 2394 1807
rect 2399 1802 2400 1807
rect 2384 1607 2400 1802
rect 2389 1602 2394 1607
rect 2399 1602 2400 1607
rect 2384 1407 2400 1602
rect 2389 1402 2394 1407
rect 2399 1402 2400 1407
rect 2384 1207 2400 1402
rect 2389 1202 2394 1207
rect 2399 1202 2400 1207
rect 2384 1007 2400 1202
rect 2389 1002 2394 1007
rect 2399 1002 2400 1007
rect 2384 807 2400 1002
rect 2389 802 2394 807
rect 2399 802 2400 807
rect 2384 607 2400 802
rect 2389 602 2394 607
rect 2399 602 2400 607
rect 2384 407 2400 602
rect 2749 452 2754 577
rect 2813 462 2818 1817
rect 2904 1707 2920 1902
rect 2909 1702 2914 1707
rect 2919 1702 2920 1707
rect 2904 1507 2920 1702
rect 3133 1572 3138 1937
rect 2909 1502 2914 1507
rect 2919 1502 2920 1507
rect 2904 1307 2920 1502
rect 2909 1302 2914 1307
rect 2919 1302 2920 1307
rect 2904 1107 2920 1302
rect 2909 1102 2914 1107
rect 2919 1102 2920 1107
rect 2877 932 2882 947
rect 2904 907 2920 1102
rect 2909 902 2914 907
rect 2919 902 2920 907
rect 2904 707 2920 902
rect 2909 702 2914 707
rect 2919 702 2920 707
rect 2904 507 2920 702
rect 2909 502 2914 507
rect 2919 502 2920 507
rect 2389 402 2394 407
rect 2399 402 2400 407
rect 2384 207 2400 402
rect 2389 202 2394 207
rect 2399 202 2400 207
rect 2384 7 2400 202
rect 2389 2 2394 7
rect 2399 2 2400 7
rect 2384 -30 2400 2
rect 2904 307 2920 502
rect 2909 302 2914 307
rect 2919 302 2920 307
rect 2904 107 2920 302
rect 3005 192 3010 1217
rect 3037 1012 3042 1097
rect 3034 1007 3042 1012
rect 3069 512 3074 1277
rect 3149 662 3154 1307
rect 3165 152 3170 697
rect 2909 102 2914 107
rect 2919 102 2920 107
rect 2904 -30 2920 102
rect 3181 82 3186 2537
rect 3408 2407 3424 2602
rect 3413 2402 3418 2407
rect 3423 2402 3424 2407
rect 3408 2207 3424 2402
rect 3413 2202 3418 2207
rect 3423 2202 3424 2207
rect 3408 2007 3424 2202
rect 3413 2002 3418 2007
rect 3423 2002 3424 2007
rect 3408 1807 3424 2002
rect 3413 1802 3418 1807
rect 3423 1802 3424 1807
rect 3325 42 3330 1387
rect 3373 1052 3378 1747
rect 3408 1607 3424 1802
rect 3413 1602 3418 1607
rect 3423 1602 3424 1607
rect 3408 1407 3424 1602
rect 3413 1402 3418 1407
rect 3423 1402 3424 1407
rect 3408 1207 3424 1402
rect 3413 1202 3418 1207
rect 3423 1202 3424 1207
rect 3389 52 3394 1137
rect 3408 1007 3424 1202
rect 3413 1002 3418 1007
rect 3423 1002 3424 1007
rect 3408 807 3424 1002
rect 3413 802 3418 807
rect 3423 802 3424 807
rect 3408 607 3424 802
rect 3437 752 3442 2027
rect 3453 1162 3458 2747
rect 3413 602 3418 607
rect 3423 602 3424 607
rect 3408 407 3424 602
rect 3413 402 3418 407
rect 3423 402 3424 407
rect 3408 207 3424 402
rect 3413 202 3418 207
rect 3423 202 3424 207
rect 3408 7 3424 202
rect 3469 72 3474 2417
rect 3501 1542 3506 3517
rect 3485 62 3490 1487
rect 3501 352 3506 1327
rect 3517 432 3522 2247
rect 3533 1552 3538 2077
rect 3565 1842 3570 3547
rect 3581 1762 3586 3087
rect 3533 1272 3538 1537
rect 3533 692 3538 1147
rect 3549 162 3554 1687
rect 3565 172 3570 1607
rect 3597 1452 3602 3437
rect 3613 1952 3618 3537
rect 3741 3462 3746 3527
rect 3581 342 3586 1117
rect 3597 352 3602 1377
rect 3613 1002 3618 1927
rect 3629 1462 3634 2367
rect 3629 1322 3634 1447
rect 3645 1382 3650 3087
rect 3661 2142 3666 3437
rect 3645 1282 3650 1357
rect 3613 742 3618 987
rect 3629 372 3634 917
rect 3645 642 3650 1257
rect 3661 362 3666 2057
rect 3677 1512 3682 2287
rect 3693 2282 3698 3077
rect 3709 2052 3714 3087
rect 3725 2542 3730 3077
rect 3677 172 3682 1487
rect 3693 1482 3698 2047
rect 3709 1642 3714 2037
rect 3677 82 3682 167
rect 3693 72 3698 1367
rect 3709 132 3714 1557
rect 3725 1332 3730 1727
rect 3725 152 3730 777
rect 3741 172 3746 1597
rect 3757 1252 3762 1937
rect 3757 72 3762 1197
rect 3773 1072 3778 1867
rect 3413 2 3418 7
rect 3423 2 3424 7
rect 3408 -30 3424 2
use BUFX2  BUFX2_62
timestamp 1719641852
transform -1 0 28 0 -1 105
box -2 -3 26 103
use DFFSR  DFFSR_91
timestamp 1719641852
transform -1 0 204 0 -1 105
box -2 -3 178 103
use BUFX2  BUFX2_68
timestamp 1719641852
transform -1 0 28 0 1 105
box -2 -3 26 103
use CLKBUF1  CLKBUF1_57
timestamp 1719641852
transform 1 0 28 0 1 105
box -2 -3 74 103
use CLKBUF1  CLKBUF1_10
timestamp 1719641852
transform -1 0 172 0 1 105
box -2 -3 74 103
use BUFX2  BUFX2_64
timestamp 1719641852
transform -1 0 196 0 1 105
box -2 -3 26 103
use CLKBUF1  CLKBUF1_20
timestamp 1719641852
transform 1 0 196 0 1 105
box -2 -3 74 103
use NAND3X1  NAND3X1_1
timestamp 1719641852
transform 1 0 252 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_76
timestamp 1719641852
transform -1 0 252 0 -1 105
box -2 -3 26 103
use BUFX2  BUFX2_67
timestamp 1719641852
transform -1 0 228 0 -1 105
box -2 -3 26 103
use CLKBUF1  CLKBUF1_60
timestamp 1719641852
transform 1 0 268 0 1 105
box -2 -3 74 103
use BUFX2  BUFX2_30
timestamp 1719641852
transform -1 0 356 0 -1 105
box -2 -3 26 103
use BUFX2  BUFX2_34
timestamp 1719641852
transform -1 0 332 0 -1 105
box -2 -3 26 103
use BUFX2  BUFX2_29
timestamp 1719641852
transform -1 0 308 0 -1 105
box -2 -3 26 103
use CLKBUF1  CLKBUF1_2
timestamp 1719641852
transform 1 0 356 0 1 105
box -2 -3 74 103
use FILL  FILL_1_0_1
timestamp 1719641852
transform 1 0 348 0 1 105
box -2 -3 10 103
use FILL  FILL_1_0_0
timestamp 1719641852
transform 1 0 340 0 1 105
box -2 -3 10 103
use FILL  FILL_0_0_1
timestamp 1719641852
transform -1 0 372 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_0_0
timestamp 1719641852
transform -1 0 364 0 -1 105
box -2 -3 10 103
use BUFX2  BUFX2_66
timestamp 1719641852
transform -1 0 396 0 -1 105
box -2 -3 26 103
use DFFSR  DFFSR_95
timestamp 1719641852
transform -1 0 572 0 -1 105
box -2 -3 178 103
use DFFSR  DFFSR_31
timestamp 1719641852
transform 1 0 428 0 1 105
box -2 -3 178 103
use BUFX2  BUFX2_27
timestamp 1719641852
transform -1 0 596 0 -1 105
box -2 -3 26 103
use BUFX2  BUFX2_32
timestamp 1719641852
transform 1 0 596 0 -1 105
box -2 -3 26 103
use BUFX2  BUFX2_51
timestamp 1719641852
transform 1 0 620 0 -1 105
box -2 -3 26 103
use DFFSR  DFFSR_80
timestamp 1719641852
transform -1 0 820 0 -1 105
box -2 -3 178 103
use OAI21X1  OAI21X1_154
timestamp 1719641852
transform 1 0 604 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_157
timestamp 1719641852
transform 1 0 636 0 1 105
box -2 -3 34 103
use BUFX2  BUFX2_33
timestamp 1719641852
transform 1 0 668 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_156
timestamp 1719641852
transform 1 0 692 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_152
timestamp 1719641852
transform 1 0 724 0 1 105
box -2 -3 34 103
use FILL  FILL_0_1_0
timestamp 1719641852
transform 1 0 820 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_1_1
timestamp 1719641852
transform 1 0 828 0 -1 105
box -2 -3 10 103
use DFFSR  DFFSR_89
timestamp 1719641852
transform 1 0 836 0 -1 105
box -2 -3 178 103
use BUFX2  BUFX2_28
timestamp 1719641852
transform 1 0 756 0 1 105
box -2 -3 26 103
use FILL  FILL_1_1_0
timestamp 1719641852
transform -1 0 788 0 1 105
box -2 -3 10 103
use FILL  FILL_1_1_1
timestamp 1719641852
transform -1 0 796 0 1 105
box -2 -3 10 103
use DFFSR  DFFSR_30
timestamp 1719641852
transform -1 0 972 0 1 105
box -2 -3 178 103
use BUFX2  BUFX2_60
timestamp 1719641852
transform 1 0 1012 0 -1 105
box -2 -3 26 103
use DFFSR  DFFSR_79
timestamp 1719641852
transform 1 0 1036 0 -1 105
box -2 -3 178 103
use OAI21X1  OAI21X1_12
timestamp 1719641852
transform 1 0 972 0 1 105
box -2 -3 34 103
use INVX1  INVX1_6
timestamp 1719641852
transform -1 0 1020 0 1 105
box -2 -3 18 103
use NAND3X1  NAND3X1_8
timestamp 1719641852
transform 1 0 1020 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_11
timestamp 1719641852
transform 1 0 1052 0 1 105
box -2 -3 34 103
use NAND3X1  NAND3X1_4
timestamp 1719641852
transform -1 0 1116 0 1 105
box -2 -3 34 103
use BUFX2  BUFX2_50
timestamp 1719641852
transform 1 0 1212 0 -1 105
box -2 -3 26 103
use DFFSR  DFFSR_94
timestamp 1719641852
transform 1 0 1236 0 -1 105
box -2 -3 178 103
use OAI21X1  OAI21X1_4
timestamp 1719641852
transform -1 0 1148 0 1 105
box -2 -3 34 103
use INVX1  INVX1_2
timestamp 1719641852
transform -1 0 1164 0 1 105
box -2 -3 18 103
use OAI21X1  OAI21X1_3
timestamp 1719641852
transform 1 0 1164 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_6
timestamp 1719641852
transform 1 0 1196 0 1 105
box -2 -3 26 103
use BUFX4  BUFX4_71
timestamp 1719641852
transform -1 0 1252 0 1 105
box -2 -3 34 103
use BUFX4  BUFX4_72
timestamp 1719641852
transform 1 0 1252 0 1 105
box -2 -3 34 103
use FILL  FILL_0_2_0
timestamp 1719641852
transform 1 0 1412 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_2_1
timestamp 1719641852
transform 1 0 1420 0 -1 105
box -2 -3 10 103
use BUFX2  BUFX2_65
timestamp 1719641852
transform 1 0 1428 0 -1 105
box -2 -3 26 103
use FILL  FILL_1_2_0
timestamp 1719641852
transform 1 0 1284 0 1 105
box -2 -3 10 103
use FILL  FILL_1_2_1
timestamp 1719641852
transform 1 0 1292 0 1 105
box -2 -3 10 103
use DFFSR  DFFSR_26
timestamp 1719641852
transform 1 0 1300 0 1 105
box -2 -3 178 103
use CLKBUF1  CLKBUF1_30
timestamp 1719641852
transform -1 0 1524 0 -1 105
box -2 -3 74 103
use BUFX2  BUFX2_61
timestamp 1719641852
transform 1 0 1524 0 -1 105
box -2 -3 26 103
use DFFSR  DFFSR_92
timestamp 1719641852
transform 1 0 1548 0 -1 105
box -2 -3 178 103
use DFFSR  DFFSR_90
timestamp 1719641852
transform -1 0 1652 0 1 105
box -2 -3 178 103
use BUFX2  BUFX2_63
timestamp 1719641852
transform 1 0 1724 0 -1 105
box -2 -3 26 103
use CLKBUF1  CLKBUF1_16
timestamp 1719641852
transform -1 0 1820 0 -1 105
box -2 -3 74 103
use DFFSR  DFFSR_206
timestamp 1719641852
transform -1 0 1828 0 1 105
box -2 -3 178 103
use FILL  FILL_0_3_0
timestamp 1719641852
transform 1 0 1820 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_3_1
timestamp 1719641852
transform 1 0 1828 0 -1 105
box -2 -3 10 103
use DFFSR  DFFSR_175
timestamp 1719641852
transform 1 0 1836 0 -1 105
box -2 -3 178 103
use CLKBUF1  CLKBUF1_33
timestamp 1719641852
transform 1 0 1828 0 1 105
box -2 -3 74 103
use FILL  FILL_1_3_0
timestamp 1719641852
transform 1 0 1900 0 1 105
box -2 -3 10 103
use FILL  FILL_1_3_1
timestamp 1719641852
transform 1 0 1908 0 1 105
box -2 -3 10 103
use DFFSR  DFFSR_177
timestamp 1719641852
transform 1 0 1916 0 1 105
box -2 -3 178 103
use DFFSR  DFFSR_178
timestamp 1719641852
transform 1 0 2012 0 -1 105
box -2 -3 178 103
use OAI21X1  OAI21X1_452
timestamp 1719641852
transform 1 0 2092 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_456
timestamp 1719641852
transform -1 0 2156 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_442
timestamp 1719641852
transform 1 0 2156 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_257
timestamp 1719641852
transform -1 0 2212 0 -1 105
box -2 -3 26 103
use DFFSR  DFFSR_207
timestamp 1719641852
transform 1 0 2212 0 -1 105
box -2 -3 178 103
use NAND2X1  NAND2X1_260
timestamp 1719641852
transform -1 0 2212 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_561
timestamp 1719641852
transform -1 0 2244 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_447
timestamp 1719641852
transform -1 0 2276 0 1 105
box -2 -3 34 103
use DFFSR  DFFSR_208
timestamp 1719641852
transform 1 0 2276 0 1 105
box -2 -3 178 103
use FILL  FILL_0_4_0
timestamp 1719641852
transform -1 0 2396 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_4_1
timestamp 1719641852
transform -1 0 2404 0 -1 105
box -2 -3 10 103
use DFFSR  DFFSR_237
timestamp 1719641852
transform -1 0 2580 0 -1 105
box -2 -3 178 103
use FILL  FILL_1_4_0
timestamp 1719641852
transform -1 0 2460 0 1 105
box -2 -3 10 103
use FILL  FILL_1_4_1
timestamp 1719641852
transform -1 0 2468 0 1 105
box -2 -3 10 103
use DFFSR  DFFSR_240
timestamp 1719641852
transform -1 0 2644 0 1 105
box -2 -3 178 103
use DFFSR  DFFSR_222
timestamp 1719641852
transform -1 0 2756 0 -1 105
box -2 -3 178 103
use NOR2X1  NOR2X1_237
timestamp 1719641852
transform 1 0 2644 0 1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_156
timestamp 1719641852
transform -1 0 2700 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_451
timestamp 1719641852
transform -1 0 2732 0 1 105
box -2 -3 34 103
use CLKBUF1  CLKBUF1_26
timestamp 1719641852
transform -1 0 2828 0 -1 105
box -2 -3 74 103
use NOR2X1  NOR2X1_233
timestamp 1719641852
transform -1 0 2852 0 -1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_232
timestamp 1719641852
transform -1 0 2876 0 -1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_151
timestamp 1719641852
transform -1 0 2908 0 -1 105
box -2 -3 34 103
use CLKBUF1  CLKBUF1_11
timestamp 1719641852
transform -1 0 2804 0 1 105
box -2 -3 74 103
use INVX8  INVX8_12
timestamp 1719641852
transform -1 0 2844 0 1 105
box -2 -3 42 103
use BUFX4  BUFX4_224
timestamp 1719641852
transform -1 0 2876 0 1 105
box -2 -3 34 103
use BUFX4  BUFX4_223
timestamp 1719641852
transform 1 0 2876 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_441
timestamp 1719641852
transform 1 0 2988 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_440
timestamp 1719641852
transform -1 0 2988 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_437
timestamp 1719641852
transform 1 0 2924 0 1 105
box -2 -3 34 103
use FILL  FILL_1_5_1
timestamp 1719641852
transform 1 0 2916 0 1 105
box -2 -3 10 103
use FILL  FILL_1_5_0
timestamp 1719641852
transform 1 0 2908 0 1 105
box -2 -3 10 103
use FILL  FILL_0_5_1
timestamp 1719641852
transform 1 0 2916 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_5_0
timestamp 1719641852
transform 1 0 2908 0 -1 105
box -2 -3 10 103
use AOI21X1  AOI21X1_153
timestamp 1719641852
transform -1 0 3052 0 1 105
box -2 -3 34 103
use DFFSR  DFFSR_224
timestamp 1719641852
transform -1 0 3228 0 1 105
box -2 -3 178 103
use DFFSR  DFFSR_210
timestamp 1719641852
transform 1 0 2924 0 -1 105
box -2 -3 178 103
use NOR2X1  NOR2X1_82
timestamp 1719641852
transform 1 0 3100 0 -1 105
box -2 -3 26 103
use INVX1  INVX1_89
timestamp 1719641852
transform -1 0 3140 0 -1 105
box -2 -3 18 103
use DFFSR  DFFSR_225
timestamp 1719641852
transform -1 0 3316 0 -1 105
box -2 -3 178 103
use CLKBUF1  CLKBUF1_56
timestamp 1719641852
transform -1 0 3300 0 1 105
box -2 -3 74 103
use NAND3X1  NAND3X1_128
timestamp 1719641852
transform -1 0 3348 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_110
timestamp 1719641852
transform 1 0 3348 0 -1 105
box -2 -3 26 103
use NAND3X1  NAND3X1_124
timestamp 1719641852
transform -1 0 3404 0 -1 105
box -2 -3 34 103
use FILL  FILL_0_6_0
timestamp 1719641852
transform -1 0 3412 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_6_1
timestamp 1719641852
transform -1 0 3420 0 -1 105
box -2 -3 10 103
use BUFX4  BUFX4_43
timestamp 1719641852
transform -1 0 3452 0 -1 105
box -2 -3 34 103
use INVX2  INVX2_152
timestamp 1719641852
transform -1 0 3316 0 1 105
box -2 -3 18 103
use DFFSR  DFFSR_209
timestamp 1719641852
transform -1 0 3492 0 1 105
box -2 -3 178 103
use NAND3X1  NAND3X1_140
timestamp 1719641852
transform -1 0 3484 0 -1 105
box -2 -3 34 103
use BUFX4  BUFX4_198
timestamp 1719641852
transform -1 0 3540 0 1 105
box -2 -3 34 103
use FILL  FILL_1_6_1
timestamp 1719641852
transform -1 0 3508 0 1 105
box -2 -3 10 103
use FILL  FILL_1_6_0
timestamp 1719641852
transform -1 0 3500 0 1 105
box -2 -3 10 103
use BUFX4  BUFX4_216
timestamp 1719641852
transform -1 0 3548 0 -1 105
box -2 -3 34 103
use BUFX4  BUFX4_186
timestamp 1719641852
transform 1 0 3484 0 -1 105
box -2 -3 34 103
use NAND3X1  NAND3X1_139
timestamp 1719641852
transform -1 0 3572 0 1 105
box -2 -3 34 103
use BUFX4  BUFX4_214
timestamp 1719641852
transform 1 0 3548 0 -1 105
box -2 -3 34 103
use BUFX4  BUFX4_46
timestamp 1719641852
transform -1 0 3604 0 1 105
box -2 -3 34 103
use INVX4  INVX4_4
timestamp 1719641852
transform 1 0 3580 0 -1 105
box -2 -3 26 103
use BUFX4  BUFX4_41
timestamp 1719641852
transform -1 0 3636 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_162
timestamp 1719641852
transform 1 0 3604 0 -1 105
box -2 -3 26 103
use BUFX4  BUFX4_44
timestamp 1719641852
transform -1 0 3668 0 1 105
box -2 -3 34 103
use BUFX4  BUFX4_184
timestamp 1719641852
transform -1 0 3684 0 -1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_68
timestamp 1719641852
transform 1 0 3628 0 -1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_29
timestamp 1719641852
transform 1 0 3668 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_204
timestamp 1719641852
transform 1 0 3684 0 -1 105
box -2 -3 34 103
use BUFX4  BUFX4_196
timestamp 1719641852
transform -1 0 3764 0 1 105
box -2 -3 34 103
use NAND3X1  NAND3X1_155
timestamp 1719641852
transform -1 0 3732 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_200
timestamp 1719641852
transform -1 0 3764 0 -1 105
box -2 -3 34 103
use INVX1  INVX1_84
timestamp 1719641852
transform -1 0 3732 0 -1 105
box -2 -3 18 103
use FILL  FILL_2_1
timestamp 1719641852
transform 1 0 3764 0 1 105
box -2 -3 10 103
use FILL  FILL_1_1
timestamp 1719641852
transform -1 0 3772 0 -1 105
box -2 -3 10 103
use FILL  FILL_2_2
timestamp 1719641852
transform 1 0 3772 0 1 105
box -2 -3 10 103
use FILL  FILL_1_2
timestamp 1719641852
transform -1 0 3780 0 -1 105
box -2 -3 10 103
use DFFSR  DFFSR_105
timestamp 1719641852
transform 1 0 4 0 -1 305
box -2 -3 178 103
use DFFSR  DFFSR_93
timestamp 1719641852
transform -1 0 356 0 -1 305
box -2 -3 178 103
use FILL  FILL_2_0_0
timestamp 1719641852
transform -1 0 364 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_0_1
timestamp 1719641852
transform -1 0 372 0 -1 305
box -2 -3 10 103
use DFFSR  DFFSR_96
timestamp 1719641852
transform -1 0 548 0 -1 305
box -2 -3 178 103
use OAI21X1  OAI21X1_153
timestamp 1719641852
transform 1 0 548 0 -1 305
box -2 -3 34 103
use CLKBUF1  CLKBUF1_8
timestamp 1719641852
transform 1 0 580 0 -1 305
box -2 -3 74 103
use OAI21X1  OAI21X1_158
timestamp 1719641852
transform -1 0 684 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_155
timestamp 1719641852
transform 1 0 684 0 -1 305
box -2 -3 34 103
use BUFX2  BUFX2_31
timestamp 1719641852
transform 1 0 716 0 -1 305
box -2 -3 26 103
use DFFSR  DFFSR_28
timestamp 1719641852
transform -1 0 916 0 -1 305
box -2 -3 178 103
use FILL  FILL_2_1_0
timestamp 1719641852
transform 1 0 916 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_1_1
timestamp 1719641852
transform 1 0 924 0 -1 305
box -2 -3 10 103
use OAI21X1  OAI21X1_8
timestamp 1719641852
transform 1 0 932 0 -1 305
box -2 -3 34 103
use INVX1  INVX1_4
timestamp 1719641852
transform -1 0 980 0 -1 305
box -2 -3 18 103
use NAND3X1  NAND3X1_6
timestamp 1719641852
transform 1 0 980 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_7
timestamp 1719641852
transform 1 0 1012 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_1
timestamp 1719641852
transform -1 0 1068 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_14
timestamp 1719641852
transform 1 0 1068 0 -1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_9
timestamp 1719641852
transform 1 0 1100 0 -1 305
box -2 -3 34 103
use INVX1  INVX1_7
timestamp 1719641852
transform 1 0 1132 0 -1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_13
timestamp 1719641852
transform 1 0 1148 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_4
timestamp 1719641852
transform 1 0 1180 0 -1 305
box -2 -3 26 103
use BUFX4  BUFX4_68
timestamp 1719641852
transform -1 0 1236 0 -1 305
box -2 -3 34 103
use DFFSR  DFFSR_145
timestamp 1719641852
transform 1 0 1236 0 -1 305
box -2 -3 178 103
use FILL  FILL_2_2_0
timestamp 1719641852
transform -1 0 1420 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_2_1
timestamp 1719641852
transform -1 0 1428 0 -1 305
box -2 -3 10 103
use MUX2X1  MUX2X1_5
timestamp 1719641852
transform -1 0 1476 0 -1 305
box -2 -3 50 103
use NAND3X1  NAND3X1_96
timestamp 1719641852
transform -1 0 1508 0 -1 305
box -2 -3 34 103
use AOI22X1  AOI22X1_21
timestamp 1719641852
transform 1 0 1508 0 -1 305
box -2 -3 42 103
use NAND3X1  NAND3X1_99
timestamp 1719641852
transform -1 0 1580 0 -1 305
box -2 -3 34 103
use AOI22X1  AOI22X1_28
timestamp 1719641852
transform -1 0 1620 0 -1 305
box -2 -3 42 103
use NAND3X1  NAND3X1_95
timestamp 1719641852
transform 1 0 1620 0 -1 305
box -2 -3 34 103
use AOI22X1  AOI22X1_20
timestamp 1719641852
transform 1 0 1652 0 -1 305
box -2 -3 42 103
use NAND3X1  NAND3X1_100
timestamp 1719641852
transform 1 0 1692 0 -1 305
box -2 -3 34 103
use AOI22X1  AOI22X1_30
timestamp 1719641852
transform 1 0 1724 0 -1 305
box -2 -3 42 103
use NAND3X1  NAND3X1_97
timestamp 1719641852
transform 1 0 1764 0 -1 305
box -2 -3 34 103
use AOI22X1  AOI22X1_24
timestamp 1719641852
transform 1 0 1796 0 -1 305
box -2 -3 42 103
use NAND2X1  NAND2X1_2
timestamp 1719641852
transform 1 0 1836 0 -1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_210
timestamp 1719641852
transform -1 0 1884 0 -1 305
box -2 -3 26 103
use FILL  FILL_2_3_0
timestamp 1719641852
transform 1 0 1884 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_3_1
timestamp 1719641852
transform 1 0 1892 0 -1 305
box -2 -3 10 103
use NAND2X1  NAND2X1_7
timestamp 1719641852
transform 1 0 1900 0 -1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_202
timestamp 1719641852
transform 1 0 1924 0 -1 305
box -2 -3 26 103
use AOI22X1  AOI22X1_19
timestamp 1719641852
transform 1 0 1948 0 -1 305
box -2 -3 42 103
use NAND2X1  NAND2X1_203
timestamp 1719641852
transform 1 0 1988 0 -1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_212
timestamp 1719641852
transform -1 0 2036 0 -1 305
box -2 -3 26 103
use INVX2  INVX2_151
timestamp 1719641852
transform 1 0 2036 0 -1 305
box -2 -3 18 103
use AOI21X1  AOI21X1_190
timestamp 1719641852
transform 1 0 2052 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_562
timestamp 1719641852
transform -1 0 2116 0 -1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_192
timestamp 1719641852
transform -1 0 2148 0 -1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_191
timestamp 1719641852
transform -1 0 2180 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_563
timestamp 1719641852
transform -1 0 2212 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_569
timestamp 1719641852
transform -1 0 2244 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_446
timestamp 1719641852
transform 1 0 2244 0 -1 305
box -2 -3 34 103
use AOI22X1  AOI22X1_23
timestamp 1719641852
transform 1 0 2276 0 -1 305
box -2 -3 42 103
use FILL  FILL_2_4_0
timestamp 1719641852
transform -1 0 2324 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_4_1
timestamp 1719641852
transform -1 0 2332 0 -1 305
box -2 -3 10 103
use DFFSR  DFFSR_176
timestamp 1719641852
transform -1 0 2508 0 -1 305
box -2 -3 178 103
use NAND2X1  NAND2X1_206
timestamp 1719641852
transform -1 0 2532 0 -1 305
box -2 -3 26 103
use AOI22X1  AOI22X1_29
timestamp 1719641852
transform 1 0 2532 0 -1 305
box -2 -3 42 103
use AOI22X1  AOI22X1_27
timestamp 1719641852
transform 1 0 2572 0 -1 305
box -2 -3 42 103
use NOR2X1  NOR2X1_240
timestamp 1719641852
transform 1 0 2612 0 -1 305
box -2 -3 26 103
use DFFSR  DFFSR_205
timestamp 1719641852
transform 1 0 2636 0 -1 305
box -2 -3 178 103
use INVX2  INVX2_143
timestamp 1719641852
transform 1 0 2812 0 -1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_331
timestamp 1719641852
transform -1 0 2860 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_449
timestamp 1719641852
transform 1 0 2860 0 -1 305
box -2 -3 34 103
use FILL  FILL_2_5_0
timestamp 1719641852
transform -1 0 2900 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_5_1
timestamp 1719641852
transform -1 0 2908 0 -1 305
box -2 -3 10 103
use OAI21X1  OAI21X1_335
timestamp 1719641852
transform -1 0 2940 0 -1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_155
timestamp 1719641852
transform -1 0 2972 0 -1 305
box -2 -3 34 103
use INVX2  INVX2_110
timestamp 1719641852
transform 1 0 2972 0 -1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_450
timestamp 1719641852
transform -1 0 3020 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_436
timestamp 1719641852
transform -1 0 3052 0 -1 305
box -2 -3 34 103
use INVX2  INVX2_66
timestamp 1719641852
transform 1 0 3052 0 -1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_439
timestamp 1719641852
transform 1 0 3068 0 -1 305
box -2 -3 34 103
use DFFSR  DFFSR_241
timestamp 1719641852
transform -1 0 3276 0 -1 305
box -2 -3 178 103
use OAI21X1  OAI21X1_435
timestamp 1719641852
transform 1 0 3276 0 -1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_150
timestamp 1719641852
transform 1 0 3308 0 -1 305
box -2 -3 34 103
use FILL  FILL_2_6_0
timestamp 1719641852
transform -1 0 3348 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_6_1
timestamp 1719641852
transform -1 0 3356 0 -1 305
box -2 -3 10 103
use DFFSR  DFFSR_242
timestamp 1719641852
transform -1 0 3532 0 -1 305
box -2 -3 178 103
use CLKBUF1  CLKBUF1_58
timestamp 1719641852
transform 1 0 3532 0 -1 305
box -2 -3 74 103
use DFFSR  DFFSR_239
timestamp 1719641852
transform -1 0 3780 0 -1 305
box -2 -3 178 103
use CLKBUF1  CLKBUF1_38
timestamp 1719641852
transform -1 0 76 0 1 305
box -2 -3 74 103
use DFFSR  DFFSR_106
timestamp 1719641852
transform 1 0 76 0 1 305
box -2 -3 178 103
use NOR2X1  NOR2X1_29
timestamp 1719641852
transform -1 0 276 0 1 305
box -2 -3 26 103
use FILL  FILL_3_0_0
timestamp 1719641852
transform 1 0 276 0 1 305
box -2 -3 10 103
use FILL  FILL_3_0_1
timestamp 1719641852
transform 1 0 284 0 1 305
box -2 -3 10 103
use DFFSR  DFFSR_104
timestamp 1719641852
transform 1 0 292 0 1 305
box -2 -3 178 103
use DFFSR  DFFSR_29
timestamp 1719641852
transform 1 0 468 0 1 305
box -2 -3 178 103
use DFFSR  DFFSR_25
timestamp 1719641852
transform -1 0 820 0 1 305
box -2 -3 178 103
use INVX1  INVX1_1
timestamp 1719641852
transform 1 0 820 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_2
timestamp 1719641852
transform 1 0 836 0 1 305
box -2 -3 34 103
use FILL  FILL_3_1_0
timestamp 1719641852
transform 1 0 868 0 1 305
box -2 -3 10 103
use FILL  FILL_3_1_1
timestamp 1719641852
transform 1 0 876 0 1 305
box -2 -3 10 103
use OAI21X1  OAI21X1_1
timestamp 1719641852
transform 1 0 884 0 1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_3
timestamp 1719641852
transform 1 0 916 0 1 305
box -2 -3 34 103
use BUFX4  BUFX4_22
timestamp 1719641852
transform 1 0 948 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_10
timestamp 1719641852
transform 1 0 980 0 1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_7
timestamp 1719641852
transform 1 0 1012 0 1 305
box -2 -3 34 103
use INVX1  INVX1_5
timestamp 1719641852
transform 1 0 1044 0 1 305
box -2 -3 18 103
use NAND3X1  NAND3X1_98
timestamp 1719641852
transform 1 0 1060 0 1 305
box -2 -3 34 103
use AOI22X1  AOI22X1_26
timestamp 1719641852
transform 1 0 1092 0 1 305
box -2 -3 42 103
use OAI21X1  OAI21X1_9
timestamp 1719641852
transform 1 0 1132 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_5
timestamp 1719641852
transform -1 0 1188 0 1 305
box -2 -3 26 103
use BUFX4  BUFX4_73
timestamp 1719641852
transform -1 0 1220 0 1 305
box -2 -3 34 103
use BUFX4  BUFX4_69
timestamp 1719641852
transform 1 0 1220 0 1 305
box -2 -3 34 103
use BUFX4  BUFX4_70
timestamp 1719641852
transform -1 0 1284 0 1 305
box -2 -3 34 103
use BUFX4  BUFX4_74
timestamp 1719641852
transform 1 0 1284 0 1 305
box -2 -3 34 103
use AOI22X1  AOI22X1_78
timestamp 1719641852
transform 1 0 1316 0 1 305
box -2 -3 42 103
use FILL  FILL_3_2_0
timestamp 1719641852
transform -1 0 1364 0 1 305
box -2 -3 10 103
use FILL  FILL_3_2_1
timestamp 1719641852
transform -1 0 1372 0 1 305
box -2 -3 10 103
use AOI21X1  AOI21X1_243
timestamp 1719641852
transform -1 0 1404 0 1 305
box -2 -3 34 103
use BUFX4  BUFX4_207
timestamp 1719641852
transform 1 0 1404 0 1 305
box -2 -3 34 103
use MUX2X1  MUX2X1_11
timestamp 1719641852
transform -1 0 1484 0 1 305
box -2 -3 50 103
use NAND2X1  NAND2X1_70
timestamp 1719641852
transform -1 0 1508 0 1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_73
timestamp 1719641852
transform 1 0 1508 0 1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_71
timestamp 1719641852
transform 1 0 1532 0 1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_69
timestamp 1719641852
transform 1 0 1556 0 1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_74
timestamp 1719641852
transform -1 0 1604 0 1 305
box -2 -3 26 103
use NOR2X1  NOR2X1_297
timestamp 1719641852
transform -1 0 1628 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_655
timestamp 1719641852
transform 1 0 1628 0 1 305
box -2 -3 34 103
use DFFSR  DFFSR_146
timestamp 1719641852
transform 1 0 1660 0 1 305
box -2 -3 178 103
use NAND2X1  NAND2X1_283
timestamp 1719641852
transform 1 0 1836 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_652
timestamp 1719641852
transform 1 0 1860 0 1 305
box -2 -3 34 103
use FILL  FILL_3_3_0
timestamp 1719641852
transform 1 0 1892 0 1 305
box -2 -3 10 103
use FILL  FILL_3_3_1
timestamp 1719641852
transform 1 0 1900 0 1 305
box -2 -3 10 103
use BUFX4  BUFX4_124
timestamp 1719641852
transform 1 0 1908 0 1 305
box -2 -3 34 103
use INVX2  INVX2_137
timestamp 1719641852
transform -1 0 1956 0 1 305
box -2 -3 18 103
use NAND2X1  NAND2X1_262
timestamp 1719641852
transform 1 0 1956 0 1 305
box -2 -3 26 103
use AOI22X1  AOI22X1_22
timestamp 1719641852
transform 1 0 1980 0 1 305
box -2 -3 42 103
use AOI22X1  AOI22X1_25
timestamp 1719641852
transform -1 0 2060 0 1 305
box -2 -3 42 103
use NOR2X1  NOR2X1_267
timestamp 1719641852
transform 1 0 2060 0 1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_204
timestamp 1719641852
transform 1 0 2084 0 1 305
box -2 -3 26 103
use NOR2X1  NOR2X1_269
timestamp 1719641852
transform 1 0 2108 0 1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_195
timestamp 1719641852
transform -1 0 2164 0 1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_194
timestamp 1719641852
transform -1 0 2196 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_565
timestamp 1719641852
transform -1 0 2228 0 1 305
box -2 -3 34 103
use INVX2  INVX2_82
timestamp 1719641852
transform -1 0 2244 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_445
timestamp 1719641852
transform -1 0 2276 0 1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_154
timestamp 1719641852
transform -1 0 2308 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_444
timestamp 1719641852
transform -1 0 2340 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_560
timestamp 1719641852
transform -1 0 2372 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_559
timestamp 1719641852
transform -1 0 2404 0 1 305
box -2 -3 34 103
use FILL  FILL_3_4_0
timestamp 1719641852
transform -1 0 2412 0 1 305
box -2 -3 10 103
use FILL  FILL_3_4_1
timestamp 1719641852
transform -1 0 2420 0 1 305
box -2 -3 10 103
use INVX2  INVX2_83
timestamp 1719641852
transform -1 0 2436 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_558
timestamp 1719641852
transform -1 0 2468 0 1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_189
timestamp 1719641852
transform -1 0 2500 0 1 305
box -2 -3 34 103
use DFFSR  DFFSR_238
timestamp 1719641852
transform -1 0 2676 0 1 305
box -2 -3 178 103
use AOI21X1  AOI21X1_159
timestamp 1719641852
transform -1 0 2708 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_333
timestamp 1719641852
transform -1 0 2740 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_348
timestamp 1719641852
transform -1 0 2772 0 1 305
box -2 -3 34 103
use INVX2  INVX2_81
timestamp 1719641852
transform 1 0 2772 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_349
timestamp 1719641852
transform 1 0 2788 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_350
timestamp 1719641852
transform 1 0 2820 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_346
timestamp 1719641852
transform -1 0 2884 0 1 305
box -2 -3 34 103
use INVX2  INVX2_141
timestamp 1719641852
transform 1 0 2884 0 1 305
box -2 -3 18 103
use FILL  FILL_3_5_0
timestamp 1719641852
transform 1 0 2900 0 1 305
box -2 -3 10 103
use FILL  FILL_3_5_1
timestamp 1719641852
transform 1 0 2908 0 1 305
box -2 -3 10 103
use OAI21X1  OAI21X1_334
timestamp 1719641852
transform 1 0 2916 0 1 305
box -2 -3 34 103
use DFFSR  DFFSR_243
timestamp 1719641852
transform 1 0 2948 0 1 305
box -2 -3 178 103
use AOI21X1  AOI21X1_152
timestamp 1719641852
transform 1 0 3124 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_328
timestamp 1719641852
transform -1 0 3188 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_329
timestamp 1719641852
transform 1 0 3188 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_330
timestamp 1719641852
transform 1 0 3220 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_326
timestamp 1719641852
transform -1 0 3284 0 1 305
box -2 -3 34 103
use INVX2  INVX2_150
timestamp 1719641852
transform 1 0 3284 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_338
timestamp 1719641852
transform -1 0 3332 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_339
timestamp 1719641852
transform -1 0 3364 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_337
timestamp 1719641852
transform -1 0 3396 0 1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_107
timestamp 1719641852
transform 1 0 3396 0 1 305
box -2 -3 34 103
use FILL  FILL_3_6_0
timestamp 1719641852
transform 1 0 3428 0 1 305
box -2 -3 10 103
use FILL  FILL_3_6_1
timestamp 1719641852
transform 1 0 3436 0 1 305
box -2 -3 10 103
use OAI21X1  OAI21X1_336
timestamp 1719641852
transform 1 0 3444 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_340
timestamp 1719641852
transform 1 0 3476 0 1 305
box -2 -3 34 103
use INVX2  INVX2_108
timestamp 1719641852
transform -1 0 3524 0 1 305
box -2 -3 18 103
use CLKBUF1  CLKBUF1_32
timestamp 1719641852
transform -1 0 3596 0 1 305
box -2 -3 74 103
use NOR2X1  NOR2X1_121
timestamp 1719641852
transform 1 0 3596 0 1 305
box -2 -3 26 103
use INVX1  INVX1_101
timestamp 1719641852
transform 1 0 3620 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_199
timestamp 1719641852
transform -1 0 3668 0 1 305
box -2 -3 34 103
use INVX8  INVX8_10
timestamp 1719641852
transform 1 0 3668 0 1 305
box -2 -3 42 103
use XNOR2X1  XNOR2X1_9
timestamp 1719641852
transform 1 0 3708 0 1 305
box -2 -3 58 103
use FILL  FILL_4_1
timestamp 1719641852
transform 1 0 3764 0 1 305
box -2 -3 10 103
use FILL  FILL_4_2
timestamp 1719641852
transform 1 0 3772 0 1 305
box -2 -3 10 103
use DFFSR  DFFSR_108
timestamp 1719641852
transform 1 0 4 0 -1 505
box -2 -3 178 103
use XNOR2X1  XNOR2X1_1
timestamp 1719641852
transform -1 0 236 0 -1 505
box -2 -3 58 103
use AND2X2  AND2X2_7
timestamp 1719641852
transform -1 0 268 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_169
timestamp 1719641852
transform -1 0 300 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_93
timestamp 1719641852
transform -1 0 324 0 -1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_94
timestamp 1719641852
transform -1 0 348 0 -1 505
box -2 -3 26 103
use FILL  FILL_4_0_0
timestamp 1719641852
transform -1 0 356 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_0_1
timestamp 1719641852
transform -1 0 364 0 -1 505
box -2 -3 10 103
use AND2X2  AND2X2_4
timestamp 1719641852
transform -1 0 396 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_80
timestamp 1719641852
transform -1 0 420 0 -1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_28
timestamp 1719641852
transform -1 0 444 0 -1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_42
timestamp 1719641852
transform -1 0 468 0 -1 505
box -2 -3 26 103
use INVX1  INVX1_72
timestamp 1719641852
transform -1 0 484 0 -1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_167
timestamp 1719641852
transform 1 0 484 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_166
timestamp 1719641852
transform 1 0 516 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_151
timestamp 1719641852
transform 1 0 548 0 -1 505
box -2 -3 34 103
use DFFSR  DFFSR_27
timestamp 1719641852
transform -1 0 756 0 -1 505
box -2 -3 178 103
use BUFX4  BUFX4_136
timestamp 1719641852
transform -1 0 788 0 -1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_5
timestamp 1719641852
transform -1 0 820 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_6
timestamp 1719641852
transform -1 0 852 0 -1 505
box -2 -3 34 103
use FILL  FILL_4_1_0
timestamp 1719641852
transform 1 0 852 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_1_1
timestamp 1719641852
transform 1 0 860 0 -1 505
box -2 -3 10 103
use INVX1  INVX1_3
timestamp 1719641852
transform 1 0 868 0 -1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_5
timestamp 1719641852
transform 1 0 884 0 -1 505
box -2 -3 34 103
use DFFSR  DFFSR_144
timestamp 1719641852
transform 1 0 916 0 -1 505
box -2 -3 178 103
use NAND2X1  NAND2X1_8
timestamp 1719641852
transform 1 0 1092 0 -1 505
box -2 -3 26 103
use AOI22X1  AOI22X1_79
timestamp 1719641852
transform -1 0 1156 0 -1 505
box -2 -3 42 103
use MUX2X1  MUX2X1_6
timestamp 1719641852
transform 1 0 1156 0 -1 505
box -2 -3 50 103
use MUX2X1  MUX2X1_7
timestamp 1719641852
transform -1 0 1252 0 -1 505
box -2 -3 50 103
use NAND3X1  NAND3X1_94
timestamp 1719641852
transform -1 0 1284 0 -1 505
box -2 -3 34 103
use BUFX4  BUFX4_21
timestamp 1719641852
transform 1 0 1284 0 -1 505
box -2 -3 34 103
use AOI22X1  AOI22X1_17
timestamp 1719641852
transform 1 0 1316 0 -1 505
box -2 -3 42 103
use INVX1  INVX1_142
timestamp 1719641852
transform -1 0 1372 0 -1 505
box -2 -3 18 103
use FILL  FILL_4_2_0
timestamp 1719641852
transform 1 0 1372 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_2_1
timestamp 1719641852
transform 1 0 1380 0 -1 505
box -2 -3 10 103
use AOI22X1  AOI22X1_32
timestamp 1719641852
transform 1 0 1388 0 -1 505
box -2 -3 42 103
use AOI22X1  AOI22X1_84
timestamp 1719641852
transform -1 0 1468 0 -1 505
box -2 -3 42 103
use NAND3X1  NAND3X1_101
timestamp 1719641852
transform -1 0 1500 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_75
timestamp 1719641852
transform -1 0 1524 0 -1 505
box -2 -3 26 103
use DFFSR  DFFSR_147
timestamp 1719641852
transform 1 0 1524 0 -1 505
box -2 -3 178 103
use INVX1  INVX1_141
timestamp 1719641852
transform -1 0 1716 0 -1 505
box -2 -3 18 103
use INVX2  INVX2_139
timestamp 1719641852
transform 1 0 1716 0 -1 505
box -2 -3 18 103
use NAND2X1  NAND2X1_201
timestamp 1719641852
transform 1 0 1732 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_660
timestamp 1719641852
transform 1 0 1756 0 -1 505
box -2 -3 34 103
use INVX1  INVX1_92
timestamp 1719641852
transform 1 0 1788 0 -1 505
box -2 -3 18 103
use AOI21X1  AOI21X1_198
timestamp 1719641852
transform 1 0 1804 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_576
timestamp 1719641852
transform 1 0 1836 0 -1 505
box -2 -3 34 103
use FILL  FILL_4_3_0
timestamp 1719641852
transform 1 0 1868 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_3_1
timestamp 1719641852
transform 1 0 1876 0 -1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_577
timestamp 1719641852
transform 1 0 1884 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_578
timestamp 1719641852
transform 1 0 1916 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_579
timestamp 1719641852
transform 1 0 1948 0 -1 505
box -2 -3 34 103
use DFFSR  DFFSR_173
timestamp 1719641852
transform -1 0 2156 0 -1 505
box -2 -3 178 103
use OAI21X1  OAI21X1_564
timestamp 1719641852
transform 1 0 2156 0 -1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_193
timestamp 1719641852
transform -1 0 2220 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_455
timestamp 1719641852
transform -1 0 2252 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_454
timestamp 1719641852
transform -1 0 2284 0 -1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_196
timestamp 1719641852
transform 1 0 2284 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_566
timestamp 1719641852
transform 1 0 2316 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_568
timestamp 1719641852
transform -1 0 2380 0 -1 505
box -2 -3 34 103
use INVX2  INVX2_69
timestamp 1719641852
transform 1 0 2380 0 -1 505
box -2 -3 18 103
use FILL  FILL_4_4_0
timestamp 1719641852
transform 1 0 2396 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_4_1
timestamp 1719641852
transform 1 0 2404 0 -1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_567
timestamp 1719641852
transform 1 0 2412 0 -1 505
box -2 -3 34 103
use INVX2  INVX2_109
timestamp 1719641852
transform 1 0 2444 0 -1 505
box -2 -3 18 103
use AOI22X1  AOI22X1_62
timestamp 1719641852
transform 1 0 2460 0 -1 505
box -2 -3 42 103
use CLKBUF1  CLKBUF1_24
timestamp 1719641852
transform 1 0 2500 0 -1 505
box -2 -3 74 103
use INVX2  INVX2_64
timestamp 1719641852
transform 1 0 2572 0 -1 505
box -2 -3 18 103
use AOI22X1  AOI22X1_69
timestamp 1719641852
transform 1 0 2588 0 -1 505
box -2 -3 42 103
use OAI21X1  OAI21X1_458
timestamp 1719641852
transform -1 0 2660 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_459
timestamp 1719641852
transform 1 0 2660 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_341
timestamp 1719641852
transform -1 0 2724 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_345
timestamp 1719641852
transform -1 0 2756 0 -1 505
box -2 -3 34 103
use BUFX4  BUFX4_138
timestamp 1719641852
transform 1 0 2756 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_318
timestamp 1719641852
transform -1 0 2820 0 -1 505
box -2 -3 34 103
use INVX2  INVX2_125
timestamp 1719641852
transform 1 0 2820 0 -1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_319
timestamp 1719641852
transform 1 0 2836 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_267
timestamp 1719641852
transform 1 0 2868 0 -1 505
box -2 -3 34 103
use FILL  FILL_4_5_0
timestamp 1719641852
transform -1 0 2908 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_5_1
timestamp 1719641852
transform -1 0 2916 0 -1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_320
timestamp 1719641852
transform -1 0 2948 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_399
timestamp 1719641852
transform -1 0 2980 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_400
timestamp 1719641852
transform 1 0 2980 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_396
timestamp 1719641852
transform -1 0 3044 0 -1 505
box -2 -3 34 103
use DFFSR  DFFSR_227
timestamp 1719641852
transform -1 0 3220 0 -1 505
box -2 -3 178 103
use OAI21X1  OAI21X1_323
timestamp 1719641852
transform -1 0 3252 0 -1 505
box -2 -3 34 103
use INVX2  INVX2_65
timestamp 1719641852
transform 1 0 3252 0 -1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_324
timestamp 1719641852
transform 1 0 3268 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_325
timestamp 1719641852
transform 1 0 3300 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_321
timestamp 1719641852
transform -1 0 3364 0 -1 505
box -2 -3 34 103
use FILL  FILL_4_6_0
timestamp 1719641852
transform 1 0 3364 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_6_1
timestamp 1719641852
transform 1 0 3372 0 -1 505
box -2 -3 10 103
use DFFSR  DFFSR_236
timestamp 1719641852
transform 1 0 3380 0 -1 505
box -2 -3 178 103
use NOR2X1  NOR2X1_119
timestamp 1719641852
transform 1 0 3556 0 -1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_81
timestamp 1719641852
transform 1 0 3580 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_211
timestamp 1719641852
transform 1 0 3604 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_237
timestamp 1719641852
transform 1 0 3636 0 -1 505
box -2 -3 34 103
use INVX1  INVX1_96
timestamp 1719641852
transform 1 0 3668 0 -1 505
box -2 -3 18 103
use NOR2X1  NOR2X1_122
timestamp 1719641852
transform 1 0 3684 0 -1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_161
timestamp 1719641852
transform -1 0 3732 0 -1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_160
timestamp 1719641852
transform -1 0 3756 0 -1 505
box -2 -3 26 103
use FILL  FILL_5_1
timestamp 1719641852
transform -1 0 3764 0 -1 505
box -2 -3 10 103
use FILL  FILL_5_2
timestamp 1719641852
transform -1 0 3772 0 -1 505
box -2 -3 10 103
use FILL  FILL_5_3
timestamp 1719641852
transform -1 0 3780 0 -1 505
box -2 -3 10 103
use DFFSR  DFFSR_114
timestamp 1719641852
transform 1 0 4 0 1 505
box -2 -3 178 103
use OAI21X1  OAI21X1_168
timestamp 1719641852
transform 1 0 180 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_170
timestamp 1719641852
transform -1 0 244 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_173
timestamp 1719641852
transform -1 0 276 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_172
timestamp 1719641852
transform -1 0 308 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_43
timestamp 1719641852
transform -1 0 332 0 1 505
box -2 -3 26 103
use INVX1  INVX1_74
timestamp 1719641852
transform 1 0 332 0 1 505
box -2 -3 18 103
use FILL  FILL_5_0_0
timestamp 1719641852
transform -1 0 356 0 1 505
box -2 -3 10 103
use FILL  FILL_5_0_1
timestamp 1719641852
transform -1 0 364 0 1 505
box -2 -3 10 103
use NAND2X1  NAND2X1_86
timestamp 1719641852
transform -1 0 388 0 1 505
box -2 -3 26 103
use NAND3X1  NAND3X1_107
timestamp 1719641852
transform 1 0 388 0 1 505
box -2 -3 34 103
use NOR3X1  NOR3X1_2
timestamp 1719641852
transform 1 0 420 0 1 505
box -2 -3 66 103
use NOR2X1  NOR2X1_41
timestamp 1719641852
transform 1 0 484 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_176
timestamp 1719641852
transform -1 0 540 0 1 505
box -2 -3 34 103
use DFFSR  DFFSR_110
timestamp 1719641852
transform -1 0 716 0 1 505
box -2 -3 178 103
use BUFX4  BUFX4_143
timestamp 1719641852
transform -1 0 748 0 1 505
box -2 -3 34 103
use CLKBUF1  CLKBUF1_28
timestamp 1719641852
transform -1 0 820 0 1 505
box -2 -3 74 103
use FILL  FILL_5_1_0
timestamp 1719641852
transform 1 0 820 0 1 505
box -2 -3 10 103
use FILL  FILL_5_1_1
timestamp 1719641852
transform 1 0 828 0 1 505
box -2 -3 10 103
use DFFSR  DFFSR_140
timestamp 1719641852
transform 1 0 836 0 1 505
box -2 -3 178 103
use NAND2X1  NAND2X1_3
timestamp 1719641852
transform -1 0 1036 0 1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_72
timestamp 1719641852
transform 1 0 1036 0 1 505
box -2 -3 26 103
use INVX1  INVX1_143
timestamp 1719641852
transform -1 0 1076 0 1 505
box -2 -3 18 103
use AOI21X1  AOI21X1_244
timestamp 1719641852
transform 1 0 1076 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_285
timestamp 1719641852
transform 1 0 1108 0 1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_68
timestamp 1719641852
transform 1 0 1132 0 1 505
box -2 -3 26 103
use AOI22X1  AOI22X1_80
timestamp 1719641852
transform 1 0 1156 0 1 505
box -2 -3 42 103
use NAND2X1  NAND2X1_286
timestamp 1719641852
transform -1 0 1220 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_245
timestamp 1719641852
transform -1 0 1252 0 1 505
box -2 -3 34 103
use INVX1  INVX1_144
timestamp 1719641852
transform -1 0 1268 0 1 505
box -2 -3 18 103
use MUX2X1  MUX2X1_8
timestamp 1719641852
transform -1 0 1316 0 1 505
box -2 -3 50 103
use BUFX4  BUFX4_127
timestamp 1719641852
transform 1 0 1316 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_284
timestamp 1719641852
transform -1 0 1372 0 1 505
box -2 -3 26 103
use FILL  FILL_5_2_0
timestamp 1719641852
transform -1 0 1380 0 1 505
box -2 -3 10 103
use FILL  FILL_5_2_1
timestamp 1719641852
transform -1 0 1388 0 1 505
box -2 -3 10 103
use AOI21X1  AOI21X1_257
timestamp 1719641852
transform -1 0 1420 0 1 505
box -2 -3 34 103
use INVX1  INVX1_162
timestamp 1719641852
transform -1 0 1436 0 1 505
box -2 -3 18 103
use NAND2X1  NAND2X1_334
timestamp 1719641852
transform -1 0 1460 0 1 505
box -2 -3 26 103
use INVX1  INVX1_148
timestamp 1719641852
transform 1 0 1460 0 1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_665
timestamp 1719641852
transform 1 0 1476 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_306
timestamp 1719641852
transform 1 0 1508 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_666
timestamp 1719641852
transform 1 0 1532 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_208
timestamp 1719641852
transform -1 0 1588 0 1 505
box -2 -3 26 103
use AOI22X1  AOI22X1_31
timestamp 1719641852
transform -1 0 1628 0 1 505
box -2 -3 42 103
use NAND2X1  NAND2X1_289
timestamp 1719641852
transform 1 0 1628 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_654
timestamp 1719641852
transform -1 0 1684 0 1 505
box -2 -3 34 103
use INVX1  INVX1_95
timestamp 1719641852
transform 1 0 1684 0 1 505
box -2 -3 18 103
use DFFSR  DFFSR_179
timestamp 1719641852
transform -1 0 1876 0 1 505
box -2 -3 178 103
use FILL  FILL_5_3_0
timestamp 1719641852
transform 1 0 1876 0 1 505
box -2 -3 10 103
use FILL  FILL_5_3_1
timestamp 1719641852
transform 1 0 1884 0 1 505
box -2 -3 10 103
use NAND2X1  NAND2X1_331
timestamp 1719641852
transform 1 0 1892 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_754
timestamp 1719641852
transform -1 0 1948 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_753
timestamp 1719641852
transform -1 0 1980 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_752
timestamp 1719641852
transform -1 0 2012 0 1 505
box -2 -3 34 103
use BUFX4  BUFX4_137
timestamp 1719641852
transform 1 0 2012 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_258
timestamp 1719641852
transform 1 0 2044 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_252
timestamp 1719641852
transform -1 0 2100 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_751
timestamp 1719641852
transform 1 0 2100 0 1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_157
timestamp 1719641852
transform 1 0 2132 0 1 505
box -2 -3 34 103
use BUFX4  BUFX4_35
timestamp 1719641852
transform 1 0 2164 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_453
timestamp 1719641852
transform 1 0 2196 0 1 505
box -2 -3 34 103
use AND2X2  AND2X2_29
timestamp 1719641852
transform 1 0 2228 0 1 505
box -2 -3 34 103
use DFFSR  DFFSR_211
timestamp 1719641852
transform -1 0 2436 0 1 505
box -2 -3 178 103
use FILL  FILL_5_4_0
timestamp 1719641852
transform -1 0 2444 0 1 505
box -2 -3 10 103
use FILL  FILL_5_4_1
timestamp 1719641852
transform -1 0 2452 0 1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_738
timestamp 1719641852
transform -1 0 2484 0 1 505
box -2 -3 34 103
use AND2X2  AND2X2_28
timestamp 1719641852
transform -1 0 2516 0 1 505
box -2 -3 34 103
use DFFSR  DFFSR_223
timestamp 1719641852
transform -1 0 2692 0 1 505
box -2 -3 178 103
use OAI21X1  OAI21X1_343
timestamp 1719641852
transform -1 0 2724 0 1 505
box -2 -3 34 103
use BUFX4  BUFX4_231
timestamp 1719641852
transform 1 0 2724 0 1 505
box -2 -3 34 103
use INVX2  INVX2_127
timestamp 1719641852
transform -1 0 2772 0 1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_344
timestamp 1719641852
transform 1 0 2772 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_249
timestamp 1719641852
transform 1 0 2804 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_108
timestamp 1719641852
transform -1 0 2860 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_342
timestamp 1719641852
transform -1 0 2892 0 1 505
box -2 -3 34 103
use FILL  FILL_5_5_0
timestamp 1719641852
transform 1 0 2892 0 1 505
box -2 -3 10 103
use FILL  FILL_5_5_1
timestamp 1719641852
transform 1 0 2900 0 1 505
box -2 -3 10 103
use AOI21X1  AOI21X1_109
timestamp 1719641852
transform 1 0 2908 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_347
timestamp 1719641852
transform -1 0 2972 0 1 505
box -2 -3 34 103
use BUFX4  BUFX4_55
timestamp 1719641852
transform -1 0 3004 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_248
timestamp 1719641852
transform 1 0 3004 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_103
timestamp 1719641852
transform 1 0 3028 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_316
timestamp 1719641852
transform 1 0 3060 0 1 505
box -2 -3 34 103
use BUFX4  BUFX4_234
timestamp 1719641852
transform -1 0 3124 0 1 505
box -2 -3 34 103
use BUFX4  BUFX4_53
timestamp 1719641852
transform 1 0 3124 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_663
timestamp 1719641852
transform -1 0 3188 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_354
timestamp 1719641852
transform 1 0 3188 0 1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_105
timestamp 1719641852
transform 1 0 3220 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_327
timestamp 1719641852
transform -1 0 3284 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_322
timestamp 1719641852
transform 1 0 3284 0 1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_104
timestamp 1719641852
transform -1 0 3348 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_355
timestamp 1719641852
transform 1 0 3348 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_351
timestamp 1719641852
transform -1 0 3412 0 1 505
box -2 -3 34 103
use FILL  FILL_5_6_0
timestamp 1719641852
transform 1 0 3412 0 1 505
box -2 -3 10 103
use FILL  FILL_5_6_1
timestamp 1719641852
transform 1 0 3420 0 1 505
box -2 -3 10 103
use NOR2X1  NOR2X1_120
timestamp 1719641852
transform 1 0 3428 0 1 505
box -2 -3 26 103
use INVX1  INVX1_120
timestamp 1719641852
transform -1 0 3468 0 1 505
box -2 -3 18 103
use NOR2X1  NOR2X1_79
timestamp 1719641852
transform -1 0 3492 0 1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_80
timestamp 1719641852
transform 1 0 3492 0 1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_139
timestamp 1719641852
transform 1 0 3516 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_210
timestamp 1719641852
transform 1 0 3540 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_236
timestamp 1719641852
transform 1 0 3572 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_114
timestamp 1719641852
transform 1 0 3604 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_141
timestamp 1719641852
transform 1 0 3636 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_99
timestamp 1719641852
transform 1 0 3668 0 1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_158
timestamp 1719641852
transform 1 0 3692 0 1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_159
timestamp 1719641852
transform 1 0 3716 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_257
timestamp 1719641852
transform 1 0 3740 0 1 505
box -2 -3 34 103
use FILL  FILL_6_1
timestamp 1719641852
transform 1 0 3772 0 1 505
box -2 -3 10 103
use DFFSR  DFFSR_113
timestamp 1719641852
transform 1 0 4 0 -1 705
box -2 -3 178 103
use NOR2X1  NOR2X1_25
timestamp 1719641852
transform -1 0 204 0 -1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_26
timestamp 1719641852
transform -1 0 228 0 -1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_79
timestamp 1719641852
transform -1 0 252 0 -1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_22
timestamp 1719641852
transform 1 0 252 0 -1 705
box -2 -3 34 103
use BUFX4  BUFX4_4
timestamp 1719641852
transform -1 0 316 0 -1 705
box -2 -3 34 103
use OR2X2  OR2X2_4
timestamp 1719641852
transform 1 0 316 0 -1 705
box -2 -3 34 103
use FILL  FILL_6_0_0
timestamp 1719641852
transform 1 0 348 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_0_1
timestamp 1719641852
transform 1 0 356 0 -1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_160
timestamp 1719641852
transform 1 0 364 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_40
timestamp 1719641852
transform -1 0 420 0 -1 705
box -2 -3 26 103
use INVX1  INVX1_71
timestamp 1719641852
transform 1 0 420 0 -1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_175
timestamp 1719641852
transform 1 0 436 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_23
timestamp 1719641852
transform 1 0 468 0 -1 705
box -2 -3 34 103
use INVX1  INVX1_75
timestamp 1719641852
transform -1 0 516 0 -1 705
box -2 -3 18 103
use INVX2  INVX2_41
timestamp 1719641852
transform -1 0 532 0 -1 705
box -2 -3 18 103
use XNOR2X1  XNOR2X1_2
timestamp 1719641852
transform -1 0 588 0 -1 705
box -2 -3 58 103
use BUFX4  BUFX4_147
timestamp 1719641852
transform 1 0 588 0 -1 705
box -2 -3 34 103
use BUFX4  BUFX4_97
timestamp 1719641852
transform -1 0 652 0 -1 705
box -2 -3 34 103
use DFFSR  DFFSR_143
timestamp 1719641852
transform 1 0 652 0 -1 705
box -2 -3 178 103
use INVX1  INVX1_8
timestamp 1719641852
transform -1 0 844 0 -1 705
box -2 -3 18 103
use FILL  FILL_6_1_0
timestamp 1719641852
transform 1 0 844 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_1_1
timestamp 1719641852
transform 1 0 852 0 -1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_15
timestamp 1719641852
transform 1 0 860 0 -1 705
box -2 -3 34 103
use DFFSR  DFFSR_141
timestamp 1719641852
transform 1 0 892 0 -1 705
box -2 -3 178 103
use DFFSR  DFFSR_142
timestamp 1719641852
transform 1 0 1068 0 -1 705
box -2 -3 178 103
use AOI22X1  AOI22X1_81
timestamp 1719641852
transform 1 0 1244 0 -1 705
box -2 -3 42 103
use AOI21X1  AOI21X1_246
timestamp 1719641852
transform -1 0 1316 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_287
timestamp 1719641852
transform -1 0 1340 0 -1 705
box -2 -3 26 103
use INVX1  INVX1_145
timestamp 1719641852
transform -1 0 1356 0 -1 705
box -2 -3 18 103
use NOR2X1  NOR2X1_300
timestamp 1719641852
transform -1 0 1380 0 -1 705
box -2 -3 26 103
use FILL  FILL_6_2_0
timestamp 1719641852
transform 1 0 1380 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_2_1
timestamp 1719641852
transform 1 0 1388 0 -1 705
box -2 -3 10 103
use NOR2X1  NOR2X1_301
timestamp 1719641852
transform 1 0 1396 0 -1 705
box -2 -3 26 103
use BUFX4  BUFX4_212
timestamp 1719641852
transform -1 0 1452 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_305
timestamp 1719641852
transform -1 0 1476 0 -1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_298
timestamp 1719641852
transform 1 0 1476 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_662
timestamp 1719641852
transform -1 0 1532 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_304
timestamp 1719641852
transform -1 0 1556 0 -1 705
box -2 -3 26 103
use INVX1  INVX1_147
timestamp 1719641852
transform -1 0 1572 0 -1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_661
timestamp 1719641852
transform -1 0 1604 0 -1 705
box -2 -3 34 103
use BUFX4  BUFX4_205
timestamp 1719641852
transform 1 0 1604 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_288
timestamp 1719641852
transform 1 0 1636 0 -1 705
box -2 -3 26 103
use DFFSR  DFFSR_174
timestamp 1719641852
transform 1 0 1660 0 -1 705
box -2 -3 178 103
use NAND2X1  NAND2X1_261
timestamp 1719641852
transform 1 0 1836 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_574
timestamp 1719641852
transform -1 0 1892 0 -1 705
box -2 -3 34 103
use FILL  FILL_6_3_0
timestamp 1719641852
transform -1 0 1900 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_3_1
timestamp 1719641852
transform -1 0 1908 0 -1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_573
timestamp 1719641852
transform -1 0 1940 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_197
timestamp 1719641852
transform 1 0 1940 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_571
timestamp 1719641852
transform 1 0 1972 0 -1 705
box -2 -3 34 103
use INVX2  INVX2_126
timestamp 1719641852
transform 1 0 2004 0 -1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_572
timestamp 1719641852
transform -1 0 2052 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_583
timestamp 1719641852
transform -1 0 2084 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_582
timestamp 1719641852
transform -1 0 2116 0 -1 705
box -2 -3 34 103
use INVX1  INVX1_138
timestamp 1719641852
transform 1 0 2116 0 -1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_581
timestamp 1719641852
transform -1 0 2164 0 -1 705
box -2 -3 34 103
use INVX2  INVX2_68
timestamp 1719641852
transform 1 0 2164 0 -1 705
box -2 -3 18 103
use CLKBUF1  CLKBUF1_42
timestamp 1719641852
transform 1 0 2180 0 -1 705
box -2 -3 74 103
use AOI22X1  AOI22X1_74
timestamp 1719641852
transform 1 0 2252 0 -1 705
box -2 -3 42 103
use OAI21X1  OAI21X1_735
timestamp 1719641852
transform 1 0 2292 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_462
timestamp 1719641852
transform -1 0 2356 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_740
timestamp 1719641852
transform -1 0 2388 0 -1 705
box -2 -3 34 103
use FILL  FILL_6_4_0
timestamp 1719641852
transform -1 0 2396 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_4_1
timestamp 1719641852
transform -1 0 2404 0 -1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_739
timestamp 1719641852
transform -1 0 2436 0 -1 705
box -2 -3 34 103
use AOI22X1  AOI22X1_73
timestamp 1719641852
transform -1 0 2476 0 -1 705
box -2 -3 42 103
use NAND2X1  NAND2X1_199
timestamp 1719641852
transform -1 0 2500 0 -1 705
box -2 -3 26 103
use BUFX4  BUFX4_38
timestamp 1719641852
transform 1 0 2500 0 -1 705
box -2 -3 34 103
use DFFSR  DFFSR_194
timestamp 1719641852
transform -1 0 2708 0 -1 705
box -2 -3 178 103
use NOR2X1  NOR2X1_258
timestamp 1719641852
transform -1 0 2732 0 -1 705
box -2 -3 26 103
use INVX2  INVX2_67
timestamp 1719641852
transform 1 0 2732 0 -1 705
box -2 -3 18 103
use AOI22X1  AOI22X1_63
timestamp 1719641852
transform -1 0 2788 0 -1 705
box -2 -3 42 103
use NAND2X1  NAND2X1_255
timestamp 1719641852
transform 1 0 2788 0 -1 705
box -2 -3 26 103
use INVX1  INVX1_133
timestamp 1719641852
transform -1 0 2828 0 -1 705
box -2 -3 18 103
use NAND2X1  NAND2X1_191
timestamp 1719641852
transform 1 0 2828 0 -1 705
box -2 -3 26 103
use AOI22X1  AOI22X1_70
timestamp 1719641852
transform -1 0 2892 0 -1 705
box -2 -3 42 103
use NAND2X1  NAND2X1_197
timestamp 1719641852
transform -1 0 2916 0 -1 705
box -2 -3 26 103
use FILL  FILL_6_5_0
timestamp 1719641852
transform 1 0 2916 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_5_1
timestamp 1719641852
transform 1 0 2924 0 -1 705
box -2 -3 10 103
use NOR2X1  NOR2X1_265
timestamp 1719641852
transform 1 0 2932 0 -1 705
box -2 -3 26 103
use INVX1  INVX1_131
timestamp 1719641852
transform 1 0 2956 0 -1 705
box -2 -3 18 103
use NAND2X1  NAND2X1_254
timestamp 1719641852
transform 1 0 2972 0 -1 705
box -2 -3 26 103
use AOI22X1  AOI22X1_59
timestamp 1719641852
transform -1 0 3036 0 -1 705
box -2 -3 42 103
use NOR2X1  NOR2X1_188
timestamp 1719641852
transform 1 0 3036 0 -1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_189
timestamp 1719641852
transform -1 0 3084 0 -1 705
box -2 -3 26 103
use AOI22X1  AOI22X1_58
timestamp 1719641852
transform 1 0 3084 0 -1 705
box -2 -3 42 103
use BUFX4  BUFX4_56
timestamp 1719641852
transform 1 0 3124 0 -1 705
box -2 -3 34 103
use AND2X2  AND2X2_22
timestamp 1719641852
transform 1 0 3156 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_353
timestamp 1719641852
transform -1 0 3220 0 -1 705
box -2 -3 34 103
use BUFX4  BUFX4_65
timestamp 1719641852
transform 1 0 3220 0 -1 705
box -2 -3 34 103
use INVX2  INVX2_165
timestamp 1719641852
transform 1 0 3252 0 -1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_352
timestamp 1719641852
transform -1 0 3300 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_110
timestamp 1719641852
transform 1 0 3300 0 -1 705
box -2 -3 34 103
use AND2X2  AND2X2_17
timestamp 1719641852
transform 1 0 3332 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_85
timestamp 1719641852
transform 1 0 3364 0 -1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_83
timestamp 1719641852
transform 1 0 3388 0 -1 705
box -2 -3 26 103
use FILL  FILL_6_6_0
timestamp 1719641852
transform 1 0 3412 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_6_1
timestamp 1719641852
transform 1 0 3420 0 -1 705
box -2 -3 10 103
use NOR2X1  NOR2X1_140
timestamp 1719641852
transform 1 0 3428 0 -1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_177
timestamp 1719641852
transform 1 0 3452 0 -1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_83
timestamp 1719641852
transform 1 0 3476 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_84
timestamp 1719641852
transform 1 0 3508 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_246
timestamp 1719641852
transform 1 0 3540 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_74
timestamp 1719641852
transform 1 0 3572 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_58
timestamp 1719641852
transform -1 0 3636 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_116
timestamp 1719641852
transform 1 0 3636 0 -1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_158
timestamp 1719641852
transform 1 0 3660 0 -1 705
box -2 -3 26 103
use AOI22X1  AOI22X1_40
timestamp 1719641852
transform 1 0 3684 0 -1 705
box -2 -3 42 103
use AOI21X1  AOI21X1_59
timestamp 1719641852
transform -1 0 3756 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_159
timestamp 1719641852
transform -1 0 3780 0 -1 705
box -2 -3 26 103
use BUFX4  BUFX4_87
timestamp 1719641852
transform -1 0 36 0 1 705
box -2 -3 34 103
use BUFX4  BUFX4_89
timestamp 1719641852
transform 1 0 36 0 1 705
box -2 -3 34 103
use AOI22X1  AOI22X1_35
timestamp 1719641852
transform 1 0 68 0 1 705
box -2 -3 42 103
use OR2X2  OR2X2_6
timestamp 1719641852
transform -1 0 140 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_25
timestamp 1719641852
transform -1 0 172 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_178
timestamp 1719641852
transform -1 0 204 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_27
timestamp 1719641852
transform 1 0 204 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_26
timestamp 1719641852
transform -1 0 268 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_171
timestamp 1719641852
transform 1 0 268 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_99
timestamp 1719641852
transform -1 0 324 0 1 705
box -2 -3 26 103
use INVX1  INVX1_76
timestamp 1719641852
transform -1 0 340 0 1 705
box -2 -3 18 103
use FILL  FILL_7_0_0
timestamp 1719641852
transform -1 0 348 0 1 705
box -2 -3 10 103
use FILL  FILL_7_0_1
timestamp 1719641852
transform -1 0 356 0 1 705
box -2 -3 10 103
use NOR2X1  NOR2X1_27
timestamp 1719641852
transform -1 0 380 0 1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_44
timestamp 1719641852
transform 1 0 380 0 1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_46
timestamp 1719641852
transform -1 0 428 0 1 705
box -2 -3 26 103
use AND2X2  AND2X2_8
timestamp 1719641852
transform -1 0 460 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_78
timestamp 1719641852
transform -1 0 484 0 1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_98
timestamp 1719641852
transform -1 0 508 0 1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_23
timestamp 1719641852
transform -1 0 532 0 1 705
box -2 -3 26 103
use DFFSR  DFFSR_109
timestamp 1719641852
transform -1 0 708 0 1 705
box -2 -3 178 103
use CLKBUF1  CLKBUF1_52
timestamp 1719641852
transform -1 0 780 0 1 705
box -2 -3 74 103
use OAI21X1  OAI21X1_16
timestamp 1719641852
transform 1 0 780 0 1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_10
timestamp 1719641852
transform 1 0 812 0 1 705
box -2 -3 34 103
use FILL  FILL_7_1_0
timestamp 1719641852
transform 1 0 844 0 1 705
box -2 -3 10 103
use FILL  FILL_7_1_1
timestamp 1719641852
transform 1 0 852 0 1 705
box -2 -3 10 103
use BUFX4  BUFX4_180
timestamp 1719641852
transform 1 0 860 0 1 705
box -2 -3 34 103
use CLKBUF1  CLKBUF1_66
timestamp 1719641852
transform -1 0 964 0 1 705
box -2 -3 74 103
use DFFSR  DFFSR_127
timestamp 1719641852
transform 1 0 964 0 1 705
box -2 -3 178 103
use NAND2X1  NAND2X1_59
timestamp 1719641852
transform -1 0 1164 0 1 705
box -2 -3 26 103
use AOI22X1  AOI22X1_82
timestamp 1719641852
transform 1 0 1164 0 1 705
box -2 -3 42 103
use NAND2X1  NAND2X1_309
timestamp 1719641852
transform -1 0 1228 0 1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_247
timestamp 1719641852
transform -1 0 1260 0 1 705
box -2 -3 34 103
use INVX1  INVX1_156
timestamp 1719641852
transform -1 0 1276 0 1 705
box -2 -3 18 103
use NOR2X1  NOR2X1_318
timestamp 1719641852
transform 1 0 1276 0 1 705
box -2 -3 26 103
use FILL  FILL_7_2_0
timestamp 1719641852
transform -1 0 1308 0 1 705
box -2 -3 10 103
use FILL  FILL_7_2_1
timestamp 1719641852
transform -1 0 1316 0 1 705
box -2 -3 10 103
use DFFSR  DFFSR_131
timestamp 1719641852
transform -1 0 1492 0 1 705
box -2 -3 178 103
use NOR2X1  NOR2X1_332
timestamp 1719641852
transform 1 0 1492 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_658
timestamp 1719641852
transform 1 0 1516 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_768
timestamp 1719641852
transform 1 0 1548 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_337
timestamp 1719641852
transform -1 0 1604 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_781
timestamp 1719641852
transform 1 0 1604 0 1 705
box -2 -3 34 103
use INVX1  INVX1_163
timestamp 1719641852
transform 1 0 1636 0 1 705
box -2 -3 18 103
use NOR2X1  NOR2X1_338
timestamp 1719641852
transform 1 0 1652 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_782
timestamp 1719641852
transform 1 0 1676 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_296
timestamp 1719641852
transform 1 0 1708 0 1 705
box -2 -3 26 103
use AOI22X1  AOI22X1_18
timestamp 1719641852
transform 1 0 1732 0 1 705
box -2 -3 42 103
use BUFX4  BUFX4_62
timestamp 1719641852
transform -1 0 1804 0 1 705
box -2 -3 34 103
use BUFX4  BUFX4_63
timestamp 1719641852
transform -1 0 1836 0 1 705
box -2 -3 34 103
use BUFX4  BUFX4_117
timestamp 1719641852
transform -1 0 1868 0 1 705
box -2 -3 34 103
use FILL  FILL_7_3_0
timestamp 1719641852
transform -1 0 1876 0 1 705
box -2 -3 10 103
use FILL  FILL_7_3_1
timestamp 1719641852
transform -1 0 1884 0 1 705
box -2 -3 10 103
use DFFSR  DFFSR_172
timestamp 1719641852
transform -1 0 2060 0 1 705
box -2 -3 178 103
use NAND2X1  NAND2X1_263
timestamp 1719641852
transform 1 0 2060 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_584
timestamp 1719641852
transform -1 0 2116 0 1 705
box -2 -3 34 103
use AND2X2  AND2X2_31
timestamp 1719641852
transform -1 0 2148 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_199
timestamp 1719641852
transform -1 0 2180 0 1 705
box -2 -3 34 103
use BUFX4  BUFX4_123
timestamp 1719641852
transform -1 0 2212 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_259
timestamp 1719641852
transform -1 0 2236 0 1 705
box -2 -3 26 103
use BUFX4  BUFX4_116
timestamp 1719641852
transform 1 0 2236 0 1 705
box -2 -3 34 103
use BUFX4  BUFX4_57
timestamp 1719641852
transform 1 0 2268 0 1 705
box -2 -3 34 103
use AND2X2  AND2X2_23
timestamp 1719641852
transform -1 0 2332 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_463
timestamp 1719641852
transform 1 0 2332 0 1 705
box -2 -3 34 103
use INVX1  INVX1_135
timestamp 1719641852
transform -1 0 2380 0 1 705
box -2 -3 18 103
use FILL  FILL_7_4_0
timestamp 1719641852
transform -1 0 2388 0 1 705
box -2 -3 10 103
use FILL  FILL_7_4_1
timestamp 1719641852
transform -1 0 2396 0 1 705
box -2 -3 10 103
use AOI21X1  AOI21X1_249
timestamp 1719641852
transform -1 0 2428 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_737
timestamp 1719641852
transform -1 0 2460 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_255
timestamp 1719641852
transform -1 0 2484 0 1 705
box -2 -3 26 103
use INVX2  INVX2_72
timestamp 1719641852
transform 1 0 2484 0 1 705
box -2 -3 18 103
use DFFSR  DFFSR_191
timestamp 1719641852
transform 1 0 2500 0 1 705
box -2 -3 178 103
use AOI21X1  AOI21X1_173
timestamp 1719641852
transform -1 0 2708 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_177
timestamp 1719641852
transform -1 0 2740 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_507
timestamp 1719641852
transform 1 0 2740 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_176
timestamp 1719641852
transform -1 0 2804 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_270
timestamp 1719641852
transform 1 0 2804 0 1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_131
timestamp 1719641852
transform 1 0 2828 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_158
timestamp 1719641852
transform -1 0 2892 0 1 705
box -2 -3 34 103
use FILL  FILL_7_5_0
timestamp 1719641852
transform -1 0 2900 0 1 705
box -2 -3 10 103
use FILL  FILL_7_5_1
timestamp 1719641852
transform -1 0 2908 0 1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_457
timestamp 1719641852
transform -1 0 2940 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_221
timestamp 1719641852
transform 1 0 2940 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_494
timestamp 1719641852
transform 1 0 2964 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_172
timestamp 1719641852
transform -1 0 3028 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_208
timestamp 1719641852
transform -1 0 3052 0 1 705
box -2 -3 26 103
use INVX1  INVX1_112
timestamp 1719641852
transform 1 0 3052 0 1 705
box -2 -3 18 103
use NOR2X1  NOR2X1_326
timestamp 1719641852
transform -1 0 3092 0 1 705
box -2 -3 26 103
use INVX2  INVX2_122
timestamp 1719641852
transform -1 0 3108 0 1 705
box -2 -3 18 103
use AOI21X1  AOI21X1_250
timestamp 1719641852
transform 1 0 3108 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_742
timestamp 1719641852
transform 1 0 3140 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_222
timestamp 1719641852
transform 1 0 3172 0 1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_132
timestamp 1719641852
transform 1 0 3196 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_397
timestamp 1719641852
transform 1 0 3228 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_204
timestamp 1719641852
transform -1 0 3284 0 1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_207
timestamp 1719641852
transform -1 0 3308 0 1 705
box -2 -3 26 103
use INVX1  INVX1_93
timestamp 1719641852
transform 1 0 3308 0 1 705
box -2 -3 18 103
use NOR2X1  NOR2X1_141
timestamp 1719641852
transform 1 0 3324 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_247
timestamp 1719641852
transform 1 0 3348 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_86
timestamp 1719641852
transform 1 0 3380 0 1 705
box -2 -3 26 103
use FILL  FILL_7_6_0
timestamp 1719641852
transform 1 0 3404 0 1 705
box -2 -3 10 103
use FILL  FILL_7_6_1
timestamp 1719641852
transform 1 0 3412 0 1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_213
timestamp 1719641852
transform 1 0 3420 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_84
timestamp 1719641852
transform 1 0 3452 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_212
timestamp 1719641852
transform 1 0 3476 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_302
timestamp 1719641852
transform 1 0 3508 0 1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_149
timestamp 1719641852
transform -1 0 3572 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_300
timestamp 1719641852
transform 1 0 3572 0 1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_117
timestamp 1719641852
transform 1 0 3604 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_115
timestamp 1719641852
transform 1 0 3636 0 1 705
box -2 -3 26 103
use NAND3X1  NAND3X1_125
timestamp 1719641852
transform -1 0 3692 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_100
timestamp 1719641852
transform 1 0 3692 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_220
timestamp 1719641852
transform 1 0 3716 0 1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_126
timestamp 1719641852
transform -1 0 3780 0 1 705
box -2 -3 34 103
use DFFSR  DFFSR_107
timestamp 1719641852
transform 1 0 4 0 -1 905
box -2 -3 178 103
use INVX1  INVX1_78
timestamp 1719641852
transform 1 0 180 0 -1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_179
timestamp 1719641852
transform 1 0 196 0 -1 905
box -2 -3 34 103
use CLKBUF1  CLKBUF1_17
timestamp 1719641852
transform -1 0 300 0 -1 905
box -2 -3 74 103
use INVX1  INVX1_73
timestamp 1719641852
transform -1 0 316 0 -1 905
box -2 -3 18 103
use BUFX4  BUFX4_2
timestamp 1719641852
transform 1 0 316 0 -1 905
box -2 -3 34 103
use FILL  FILL_8_0_0
timestamp 1719641852
transform 1 0 348 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_0_1
timestamp 1719641852
transform 1 0 356 0 -1 905
box -2 -3 10 103
use NOR2X1  NOR2X1_45
timestamp 1719641852
transform 1 0 364 0 -1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_21
timestamp 1719641852
transform 1 0 388 0 -1 905
box -2 -3 34 103
use AOI22X1  AOI22X1_34
timestamp 1719641852
transform -1 0 460 0 -1 905
box -2 -3 42 103
use NOR2X1  NOR2X1_24
timestamp 1719641852
transform 1 0 460 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_177
timestamp 1719641852
transform -1 0 516 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_24
timestamp 1719641852
transform 1 0 516 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_174
timestamp 1719641852
transform 1 0 548 0 -1 905
box -2 -3 34 103
use CLKBUF1  CLKBUF1_14
timestamp 1719641852
transform -1 0 652 0 -1 905
box -2 -3 74 103
use DFFSR  DFFSR_32
timestamp 1719641852
transform -1 0 828 0 -1 905
box -2 -3 178 103
use FILL  FILL_8_1_0
timestamp 1719641852
transform 1 0 828 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_1_1
timestamp 1719641852
transform 1 0 836 0 -1 905
box -2 -3 10 103
use CLKBUF1  CLKBUF1_34
timestamp 1719641852
transform 1 0 844 0 -1 905
box -2 -3 74 103
use DFFSR  DFFSR_158
timestamp 1719641852
transform -1 0 1092 0 -1 905
box -2 -3 178 103
use MUX2X1  MUX2X1_9
timestamp 1719641852
transform -1 0 1140 0 -1 905
box -2 -3 50 103
use AOI21X1  AOI21X1_18
timestamp 1719641852
transform -1 0 1172 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_310
timestamp 1719641852
transform -1 0 1196 0 -1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_16
timestamp 1719641852
transform -1 0 1228 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_58
timestamp 1719641852
transform 1 0 1228 0 -1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_15
timestamp 1719641852
transform -1 0 1284 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_319
timestamp 1719641852
transform 1 0 1284 0 -1 905
box -2 -3 26 103
use FILL  FILL_8_2_0
timestamp 1719641852
transform -1 0 1316 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_2_1
timestamp 1719641852
transform -1 0 1324 0 -1 905
box -2 -3 10 103
use DFFSR  DFFSR_130
timestamp 1719641852
transform -1 0 1500 0 -1 905
box -2 -3 178 103
use OAI21X1  OAI21X1_659
timestamp 1719641852
transform 1 0 1500 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_622
timestamp 1719641852
transform -1 0 1564 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_274
timestamp 1719641852
transform -1 0 1588 0 -1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_225
timestamp 1719641852
transform 1 0 1588 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_286
timestamp 1719641852
transform -1 0 1644 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_695
timestamp 1719641852
transform -1 0 1676 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_315
timestamp 1719641852
transform -1 0 1700 0 -1 905
box -2 -3 26 103
use INVX1  INVX1_154
timestamp 1719641852
transform -1 0 1716 0 -1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_694
timestamp 1719641852
transform -1 0 1748 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_314
timestamp 1719641852
transform -1 0 1772 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_653
timestamp 1719641852
transform 1 0 1772 0 -1 905
box -2 -3 34 103
use BUFX4  BUFX4_131
timestamp 1719641852
transform -1 0 1836 0 -1 905
box -2 -3 34 103
use AOI22X1  AOI22X1_75
timestamp 1719641852
transform 1 0 1836 0 -1 905
box -2 -3 42 103
use FILL  FILL_8_3_0
timestamp 1719641852
transform -1 0 1884 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_3_1
timestamp 1719641852
transform -1 0 1892 0 -1 905
box -2 -3 10 103
use INVX1  INVX1_139
timestamp 1719641852
transform -1 0 1908 0 -1 905
box -2 -3 18 103
use AOI22X1  AOI22X1_60
timestamp 1719641852
transform -1 0 1948 0 -1 905
box -2 -3 42 103
use DFFSR  DFFSR_190
timestamp 1719641852
transform -1 0 2124 0 -1 905
box -2 -3 178 103
use DFFSR  DFFSR_204
timestamp 1719641852
transform -1 0 2300 0 -1 905
box -2 -3 178 103
use OAI21X1  OAI21X1_460
timestamp 1719641852
transform 1 0 2300 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_464
timestamp 1719641852
transform -1 0 2364 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_273
timestamp 1719641852
transform 1 0 2364 0 -1 905
box -2 -3 26 103
use FILL  FILL_8_4_0
timestamp 1719641852
transform -1 0 2396 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_4_1
timestamp 1719641852
transform -1 0 2404 0 -1 905
box -2 -3 10 103
use OAI21X1  OAI21X1_461
timestamp 1719641852
transform -1 0 2436 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_160
timestamp 1719641852
transform -1 0 2468 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_325
timestamp 1719641852
transform 1 0 2468 0 -1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_328
timestamp 1719641852
transform -1 0 2516 0 -1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_236
timestamp 1719641852
transform 1 0 2516 0 -1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_268
timestamp 1719641852
transform 1 0 2540 0 -1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_259
timestamp 1719641852
transform 1 0 2564 0 -1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_179
timestamp 1719641852
transform -1 0 2620 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_510
timestamp 1719641852
transform 1 0 2620 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_178
timestamp 1719641852
transform 1 0 2652 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_512
timestamp 1719641852
transform 1 0 2684 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_509
timestamp 1719641852
transform -1 0 2748 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_200
timestamp 1719641852
transform 1 0 2748 0 -1 905
box -2 -3 26 103
use AOI22X1  AOI22X1_76
timestamp 1719641852
transform 1 0 2772 0 -1 905
box -2 -3 42 103
use OAI21X1  OAI21X1_448
timestamp 1719641852
transform 1 0 2812 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_394
timestamp 1719641852
transform 1 0 2844 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_129
timestamp 1719641852
transform -1 0 2908 0 -1 905
box -2 -3 34 103
use FILL  FILL_8_5_0
timestamp 1719641852
transform 1 0 2908 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_5_1
timestamp 1719641852
transform 1 0 2916 0 -1 905
box -2 -3 10 103
use NOR2X1  NOR2X1_238
timestamp 1719641852
transform 1 0 2924 0 -1 905
box -2 -3 26 103
use INVX2  INVX2_111
timestamp 1719641852
transform 1 0 2948 0 -1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_434
timestamp 1719641852
transform -1 0 2996 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_234
timestamp 1719641852
transform -1 0 3020 0 -1 905
box -2 -3 26 103
use INVX2  INVX2_70
timestamp 1719641852
transform 1 0 3020 0 -1 905
box -2 -3 18 103
use OR2X2  OR2X2_14
timestamp 1719641852
transform 1 0 3036 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_744
timestamp 1719641852
transform -1 0 3100 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_741
timestamp 1719641852
transform -1 0 3132 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_745
timestamp 1719641852
transform 1 0 3132 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_384
timestamp 1719641852
transform 1 0 3164 0 -1 905
box -2 -3 34 103
use INVX1  INVX1_130
timestamp 1719641852
transform -1 0 3212 0 -1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_388
timestamp 1719641852
transform -1 0 3244 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_127
timestamp 1719641852
transform 1 0 3244 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_210
timestamp 1719641852
transform 1 0 3276 0 -1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_137
timestamp 1719641852
transform 1 0 3300 0 -1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_138
timestamp 1719641852
transform 1 0 3324 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_245
timestamp 1719641852
transform 1 0 3348 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_125
timestamp 1719641852
transform 1 0 3380 0 -1 905
box -2 -3 26 103
use INVX1  INVX1_97
timestamp 1719641852
transform 1 0 3404 0 -1 905
box -2 -3 18 103
use FILL  FILL_8_6_0
timestamp 1719641852
transform 1 0 3420 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_6_1
timestamp 1719641852
transform 1 0 3428 0 -1 905
box -2 -3 10 103
use NOR2X1  NOR2X1_126
timestamp 1719641852
transform 1 0 3436 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_239
timestamp 1719641852
transform 1 0 3460 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_301
timestamp 1719641852
transform -1 0 3524 0 -1 905
box -2 -3 34 103
use INVX1  INVX1_94
timestamp 1719641852
transform 1 0 3524 0 -1 905
box -2 -3 18 103
use NOR2X1  NOR2X1_90
timestamp 1719641852
transform 1 0 3540 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_215
timestamp 1719641852
transform 1 0 3564 0 -1 905
box -2 -3 34 103
use BUFX4  BUFX4_218
timestamp 1719641852
transform -1 0 3628 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_227
timestamp 1719641852
transform 1 0 3628 0 -1 905
box -2 -3 34 103
use BUFX4  BUFX4_40
timestamp 1719641852
transform -1 0 3692 0 -1 905
box -2 -3 34 103
use AND2X2  AND2X2_13
timestamp 1719641852
transform 1 0 3692 0 -1 905
box -2 -3 34 103
use BUFX4  BUFX4_187
timestamp 1719641852
transform -1 0 3756 0 -1 905
box -2 -3 34 103
use FILL  FILL_9_1
timestamp 1719641852
transform -1 0 3764 0 -1 905
box -2 -3 10 103
use FILL  FILL_9_2
timestamp 1719641852
transform -1 0 3772 0 -1 905
box -2 -3 10 103
use FILL  FILL_9_3
timestamp 1719641852
transform -1 0 3780 0 -1 905
box -2 -3 10 103
use BUFX4  BUFX4_90
timestamp 1719641852
transform -1 0 36 0 1 905
box -2 -3 34 103
use DFFSR  DFFSR_111
timestamp 1719641852
transform 1 0 36 0 1 905
box -2 -3 178 103
use INVX1  INVX1_77
timestamp 1719641852
transform 1 0 212 0 1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_180
timestamp 1719641852
transform 1 0 228 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_95
timestamp 1719641852
transform 1 0 260 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_96
timestamp 1719641852
transform -1 0 308 0 1 905
box -2 -3 26 103
use BUFX4  BUFX4_3
timestamp 1719641852
transform 1 0 308 0 1 905
box -2 -3 34 103
use FILL  FILL_9_0_0
timestamp 1719641852
transform 1 0 340 0 1 905
box -2 -3 10 103
use FILL  FILL_9_0_1
timestamp 1719641852
transform 1 0 348 0 1 905
box -2 -3 10 103
use BUFX4  BUFX4_1
timestamp 1719641852
transform 1 0 356 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_31
timestamp 1719641852
transform -1 0 412 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_81
timestamp 1719641852
transform -1 0 436 0 1 905
box -2 -3 26 103
use NAND3X1  NAND3X1_106
timestamp 1719641852
transform -1 0 468 0 1 905
box -2 -3 34 103
use AOI22X1  AOI22X1_33
timestamp 1719641852
transform 1 0 468 0 1 905
box -2 -3 42 103
use OR2X2  OR2X2_5
timestamp 1719641852
transform -1 0 540 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_97
timestamp 1719641852
transform -1 0 564 0 1 905
box -2 -3 26 103
use DFFSR  DFFSR_61
timestamp 1719641852
transform -1 0 740 0 1 905
box -2 -3 178 103
use DFFSR  DFFSR_16
timestamp 1719641852
transform 1 0 740 0 1 905
box -2 -3 178 103
use FILL  FILL_9_1_0
timestamp 1719641852
transform -1 0 924 0 1 905
box -2 -3 10 103
use FILL  FILL_9_1_1
timestamp 1719641852
transform -1 0 932 0 1 905
box -2 -3 10 103
use OAI21X1  OAI21X1_48
timestamp 1719641852
transform -1 0 964 0 1 905
box -2 -3 34 103
use DFFSR  DFFSR_126
timestamp 1719641852
transform 1 0 964 0 1 905
box -2 -3 178 103
use AOI22X1  AOI22X1_83
timestamp 1719641852
transform 1 0 1140 0 1 905
box -2 -3 42 103
use AOI21X1  AOI21X1_248
timestamp 1719641852
transform -1 0 1212 0 1 905
box -2 -3 34 103
use INVX1  INVX1_157
timestamp 1719641852
transform -1 0 1228 0 1 905
box -2 -3 18 103
use DFFSR  DFFSR_124
timestamp 1719641852
transform -1 0 1404 0 1 905
box -2 -3 178 103
use FILL  FILL_9_2_0
timestamp 1719641852
transform 1 0 1404 0 1 905
box -2 -3 10 103
use FILL  FILL_9_2_1
timestamp 1719641852
transform 1 0 1412 0 1 905
box -2 -3 10 103
use NOR2X1  NOR2X1_299
timestamp 1719641852
transform 1 0 1420 0 1 905
box -2 -3 26 103
use INVX1  INVX1_60
timestamp 1719641852
transform -1 0 1460 0 1 905
box -2 -3 18 103
use CLKBUF1  CLKBUF1_45
timestamp 1719641852
transform -1 0 1532 0 1 905
box -2 -3 74 103
use AOI21X1  AOI21X1_223
timestamp 1719641852
transform -1 0 1564 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_656
timestamp 1719641852
transform 1 0 1564 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_224
timestamp 1719641852
transform 1 0 1596 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_623
timestamp 1719641852
transform -1 0 1660 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_306
timestamp 1719641852
transform 1 0 1660 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_337
timestamp 1719641852
transform 1 0 1684 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_780
timestamp 1719641852
transform -1 0 1740 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_34
timestamp 1719641852
transform 1 0 1740 0 1 905
box -2 -3 34 103
use INVX2  INVX2_71
timestamp 1719641852
transform -1 0 1788 0 1 905
box -2 -3 18 103
use INVX1  INVX1_50
timestamp 1719641852
transform -1 0 1804 0 1 905
box -2 -3 18 103
use INVX1  INVX1_98
timestamp 1719641852
transform -1 0 1820 0 1 905
box -2 -3 18 103
use AOI22X1  AOI22X1_71
timestamp 1719641852
transform -1 0 1860 0 1 905
box -2 -3 42 103
use NOR2X1  NOR2X1_272
timestamp 1719641852
transform 1 0 1860 0 1 905
box -2 -3 26 103
use FILL  FILL_9_3_0
timestamp 1719641852
transform 1 0 1884 0 1 905
box -2 -3 10 103
use FILL  FILL_9_3_1
timestamp 1719641852
transform 1 0 1892 0 1 905
box -2 -3 10 103
use OAI21X1  OAI21X1_570
timestamp 1719641852
transform 1 0 1900 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_271
timestamp 1719641852
transform -1 0 1956 0 1 905
box -2 -3 26 103
use BUFX4  BUFX4_29
timestamp 1719641852
transform 1 0 1956 0 1 905
box -2 -3 34 103
use DFFSR  DFFSR_195
timestamp 1719641852
transform 1 0 1988 0 1 905
box -2 -3 178 103
use AOI22X1  AOI22X1_61
timestamp 1719641852
transform 1 0 2164 0 1 905
box -2 -3 42 103
use NAND2X1  NAND2X1_190
timestamp 1719641852
transform 1 0 2204 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_198
timestamp 1719641852
transform 1 0 2228 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_755
timestamp 1719641852
transform 1 0 2252 0 1 905
box -2 -3 34 103
use INVX2  INVX2_124
timestamp 1719641852
transform 1 0 2284 0 1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_759
timestamp 1719641852
transform -1 0 2332 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_758
timestamp 1719641852
transform -1 0 2364 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_757
timestamp 1719641852
transform -1 0 2396 0 1 905
box -2 -3 34 103
use FILL  FILL_9_4_0
timestamp 1719641852
transform 1 0 2396 0 1 905
box -2 -3 10 103
use FILL  FILL_9_4_1
timestamp 1719641852
transform 1 0 2404 0 1 905
box -2 -3 10 103
use BUFX4  BUFX4_168
timestamp 1719641852
transform 1 0 2412 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_253
timestamp 1719641852
transform -1 0 2476 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_756
timestamp 1719641852
transform -1 0 2508 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_266
timestamp 1719641852
transform 1 0 2508 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_511
timestamp 1719641852
transform 1 0 2532 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_395
timestamp 1719641852
transform -1 0 2596 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_130
timestamp 1719641852
transform 1 0 2596 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_174
timestamp 1719641852
transform -1 0 2652 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_256
timestamp 1719641852
transform -1 0 2676 0 1 905
box -2 -3 26 103
use INVX2  INVX2_63
timestamp 1719641852
transform -1 0 2692 0 1 905
box -2 -3 18 103
use BUFX4  BUFX4_229
timestamp 1719641852
transform -1 0 2724 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_508
timestamp 1719641852
transform -1 0 2756 0 1 905
box -2 -3 34 103
use INVX2  INVX2_113
timestamp 1719641852
transform 1 0 2756 0 1 905
box -2 -3 18 103
use AOI22X1  AOI22X1_64
timestamp 1719641852
transform 1 0 2772 0 1 905
box -2 -3 42 103
use NAND2X1  NAND2X1_192
timestamp 1719641852
transform 1 0 2812 0 1 905
box -2 -3 26 103
use AOI22X1  AOI22X1_65
timestamp 1719641852
transform -1 0 2876 0 1 905
box -2 -3 42 103
use OAI21X1  OAI21X1_315
timestamp 1719641852
transform 1 0 2876 0 1 905
box -2 -3 34 103
use FILL  FILL_9_5_0
timestamp 1719641852
transform 1 0 2908 0 1 905
box -2 -3 10 103
use FILL  FILL_9_5_1
timestamp 1719641852
transform 1 0 2916 0 1 905
box -2 -3 10 103
use OAI21X1  OAI21X1_309
timestamp 1719641852
transform 1 0 2924 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_398
timestamp 1719641852
transform -1 0 2988 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_314
timestamp 1719641852
transform 1 0 2988 0 1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_209
timestamp 1719641852
transform 1 0 3020 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_308
timestamp 1719641852
transform 1 0 3052 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_106
timestamp 1719641852
transform 1 0 3084 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_332
timestamp 1719641852
transform 1 0 3116 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_207
timestamp 1719641852
transform -1 0 3172 0 1 905
box -2 -3 26 103
use INVX2  INVX2_153
timestamp 1719641852
transform -1 0 3188 0 1 905
box -2 -3 18 103
use NAND2X1  NAND2X1_205
timestamp 1719641852
transform 1 0 3188 0 1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_219
timestamp 1719641852
transform 1 0 3212 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_385
timestamp 1719641852
transform 1 0 3236 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_87
timestamp 1719641852
transform 1 0 3268 0 1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_123
timestamp 1719641852
transform 1 0 3292 0 1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_124
timestamp 1719641852
transform 1 0 3316 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_238
timestamp 1719641852
transform 1 0 3340 0 1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_148
timestamp 1719641852
transform -1 0 3404 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_88
timestamp 1719641852
transform -1 0 3428 0 1 905
box -2 -3 26 103
use FILL  FILL_9_6_0
timestamp 1719641852
transform 1 0 3428 0 1 905
box -2 -3 10 103
use FILL  FILL_9_6_1
timestamp 1719641852
transform 1 0 3436 0 1 905
box -2 -3 10 103
use OAI21X1  OAI21X1_214
timestamp 1719641852
transform 1 0 3444 0 1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_142
timestamp 1719641852
transform -1 0 3508 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_89
timestamp 1719641852
transform 1 0 3508 0 1 905
box -2 -3 26 103
use NAND3X1  NAND3X1_150
timestamp 1719641852
transform -1 0 3564 0 1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_118
timestamp 1719641852
transform -1 0 3596 0 1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_119
timestamp 1719641852
transform -1 0 3628 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_117
timestamp 1719641852
transform 1 0 3628 0 1 905
box -2 -3 26 103
use NAND3X1  NAND3X1_143
timestamp 1719641852
transform -1 0 3684 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_228
timestamp 1719641852
transform 1 0 3684 0 1 905
box -2 -3 34 103
use AND2X2  AND2X2_14
timestamp 1719641852
transform 1 0 3716 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_229
timestamp 1719641852
transform 1 0 3748 0 1 905
box -2 -3 34 103
use BUFX2  BUFX2_18
timestamp 1719641852
transform -1 0 28 0 -1 1105
box -2 -3 26 103
use BUFX2  BUFX2_13
timestamp 1719641852
transform -1 0 52 0 -1 1105
box -2 -3 26 103
use DFFSR  DFFSR_115
timestamp 1719641852
transform 1 0 52 0 -1 1105
box -2 -3 178 103
use NAND2X1  NAND2X1_84
timestamp 1719641852
transform 1 0 228 0 -1 1105
box -2 -3 26 103
use AND2X2  AND2X2_5
timestamp 1719641852
transform 1 0 252 0 -1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_102
timestamp 1719641852
transform -1 0 316 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_65
timestamp 1719641852
transform -1 0 332 0 -1 1105
box -2 -3 18 103
use FILL  FILL_10_0_0
timestamp 1719641852
transform -1 0 340 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_0_1
timestamp 1719641852
transform -1 0 348 0 -1 1105
box -2 -3 10 103
use DFFSR  DFFSR_100
timestamp 1719641852
transform -1 0 524 0 -1 1105
box -2 -3 178 103
use DFFSR  DFFSR_112
timestamp 1719641852
transform -1 0 700 0 -1 1105
box -2 -3 178 103
use OAI21X1  OAI21X1_137
timestamp 1719641852
transform 1 0 700 0 -1 1105
box -2 -3 34 103
use DFFSR  DFFSR_11
timestamp 1719641852
transform -1 0 908 0 -1 1105
box -2 -3 178 103
use FILL  FILL_10_1_0
timestamp 1719641852
transform -1 0 916 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_1_1
timestamp 1719641852
transform -1 0 924 0 -1 1105
box -2 -3 10 103
use NAND3X1  NAND3X1_26
timestamp 1719641852
transform -1 0 956 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_142
timestamp 1719641852
transform -1 0 988 0 -1 1105
box -2 -3 34 103
use INVX2  INVX2_8
timestamp 1719641852
transform 1 0 988 0 -1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_47
timestamp 1719641852
transform -1 0 1036 0 -1 1105
box -2 -3 34 103
use CLKBUF1  CLKBUF1_43
timestamp 1719641852
transform -1 0 1108 0 -1 1105
box -2 -3 74 103
use OAI22X1  OAI22X1_38
timestamp 1719641852
transform 1 0 1108 0 -1 1105
box -2 -3 42 103
use BUFX4  BUFX4_133
timestamp 1719641852
transform 1 0 1148 0 -1 1105
box -2 -3 34 103
use MUX2X1  MUX2X1_10
timestamp 1719641852
transform -1 0 1228 0 -1 1105
box -2 -3 50 103
use OAI22X1  OAI22X1_35
timestamp 1719641852
transform 1 0 1228 0 -1 1105
box -2 -3 42 103
use CLKBUF1  CLKBUF1_31
timestamp 1719641852
transform -1 0 1340 0 -1 1105
box -2 -3 74 103
use NAND2X1  NAND2X1_235
timestamp 1719641852
transform 1 0 1340 0 -1 1105
box -2 -3 26 103
use FILL  FILL_10_2_0
timestamp 1719641852
transform -1 0 1372 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_2_1
timestamp 1719641852
transform -1 0 1380 0 -1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_710
timestamp 1719641852
transform -1 0 1412 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_709
timestamp 1719641852
transform -1 0 1444 0 -1 1105
box -2 -3 34 103
use OR2X2  OR2X2_19
timestamp 1719641852
transform -1 0 1476 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_708
timestamp 1719641852
transform -1 0 1508 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_316
timestamp 1719641852
transform -1 0 1532 0 -1 1105
box -2 -3 26 103
use BUFX4  BUFX4_210
timestamp 1719641852
transform 1 0 1532 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_259
timestamp 1719641852
transform -1 0 1596 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_271
timestamp 1719641852
transform -1 0 1620 0 -1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_335
timestamp 1719641852
transform 1 0 1620 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_770
timestamp 1719641852
transform -1 0 1676 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_657
timestamp 1719641852
transform 1 0 1676 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_664
timestamp 1719641852
transform 1 0 1708 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_283
timestamp 1719641852
transform -1 0 1764 0 -1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_215
timestamp 1719641852
transform -1 0 1796 0 -1 1105
box -2 -3 34 103
use FILL  FILL_10_3_0
timestamp 1719641852
transform 1 0 1796 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_3_1
timestamp 1719641852
transform 1 0 1804 0 -1 1105
box -2 -3 10 103
use DFFSR  DFFSR_162
timestamp 1719641852
transform 1 0 1812 0 -1 1105
box -2 -3 178 103
use INVX2  INVX2_61
timestamp 1719641852
transform 1 0 1988 0 -1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_612
timestamp 1719641852
transform 1 0 2004 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_693
timestamp 1719641852
transform -1 0 2068 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_213
timestamp 1719641852
transform -1 0 2100 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_270
timestamp 1719641852
transform -1 0 2124 0 -1 1105
box -2 -3 26 103
use INVX1  INVX1_63
timestamp 1719641852
transform -1 0 2140 0 -1 1105
box -2 -3 18 103
use INVX1  INVX1_140
timestamp 1719641852
transform -1 0 2156 0 -1 1105
box -2 -3 18 103
use NOR2X1  NOR2X1_273
timestamp 1719641852
transform 1 0 2156 0 -1 1105
box -2 -3 26 103
use INVX1  INVX1_91
timestamp 1719641852
transform -1 0 2196 0 -1 1105
box -2 -3 18 103
use BUFX4  BUFX4_118
timestamp 1719641852
transform 1 0 2196 0 -1 1105
box -2 -3 34 103
use AOI22X1  AOI22X1_72
timestamp 1719641852
transform -1 0 2268 0 -1 1105
box -2 -3 42 103
use NOR2X1  NOR2X1_285
timestamp 1719641852
transform -1 0 2292 0 -1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_222
timestamp 1719641852
transform -1 0 2324 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_221
timestamp 1719641852
transform -1 0 2356 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_620
timestamp 1719641852
transform 1 0 2356 0 -1 1105
box -2 -3 34 103
use FILL  FILL_10_4_0
timestamp 1719641852
transform -1 0 2396 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_4_1
timestamp 1719641852
transform -1 0 2404 0 -1 1105
box -2 -3 10 103
use AOI21X1  AOI21X1_220
timestamp 1719641852
transform -1 0 2436 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_621
timestamp 1719641852
transform -1 0 2468 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_521
timestamp 1719641852
transform -1 0 2500 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_242
timestamp 1719641852
transform 1 0 2500 0 -1 1105
box -2 -3 26 103
use AND2X2  AND2X2_30
timestamp 1719641852
transform -1 0 2556 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_329
timestamp 1719641852
transform 1 0 2556 0 -1 1105
box -2 -3 26 103
use INVX2  INVX2_62
timestamp 1719641852
transform 1 0 2580 0 -1 1105
box -2 -3 18 103
use INVX1  INVX1_134
timestamp 1719641852
transform -1 0 2612 0 -1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_580
timestamp 1719641852
transform -1 0 2644 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_495
timestamp 1719641852
transform -1 0 2676 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_496
timestamp 1719641852
transform 1 0 2676 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_736
timestamp 1719641852
transform 1 0 2708 0 -1 1105
box -2 -3 34 103
use INVX2  INVX2_112
timestamp 1719641852
transform 1 0 2740 0 -1 1105
box -2 -3 18 103
use NOR2X1  NOR2X1_241
timestamp 1719641852
transform 1 0 2756 0 -1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_124
timestamp 1719641852
transform -1 0 2812 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_382
timestamp 1719641852
transform -1 0 2844 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_230
timestamp 1719641852
transform 1 0 2844 0 -1 1105
box -2 -3 26 103
use BUFX4  BUFX4_222
timestamp 1719641852
transform -1 0 2900 0 -1 1105
box -2 -3 34 103
use FILL  FILL_10_5_0
timestamp 1719641852
transform -1 0 2908 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_5_1
timestamp 1719641852
transform -1 0 2916 0 -1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_743
timestamp 1719641852
transform -1 0 2948 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_209
timestamp 1719641852
transform -1 0 2972 0 -1 1105
box -2 -3 26 103
use BUFX4  BUFX4_240
timestamp 1719641852
transform 1 0 2972 0 -1 1105
box -2 -3 34 103
use BUFX4  BUFX4_233
timestamp 1719641852
transform 1 0 3004 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_187
timestamp 1719641852
transform 1 0 3036 0 -1 1105
box -2 -3 26 103
use INVX1  INVX1_111
timestamp 1719641852
transform -1 0 3076 0 -1 1105
box -2 -3 18 103
use NAND3X1  NAND3X1_206
timestamp 1719641852
transform 1 0 3076 0 -1 1105
box -2 -3 34 103
use AOI22X1  AOI22X1_77
timestamp 1719641852
transform -1 0 3148 0 -1 1105
box -2 -3 42 103
use BUFX4  BUFX4_242
timestamp 1719641852
transform 1 0 3148 0 -1 1105
box -2 -3 34 103
use MUX2X1  MUX2X1_3
timestamp 1719641852
transform -1 0 3228 0 -1 1105
box -2 -3 50 103
use AOI21X1  AOI21X1_65
timestamp 1719641852
transform 1 0 3228 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_168
timestamp 1719641852
transform 1 0 3260 0 -1 1105
box -2 -3 26 103
use MUX2X1  MUX2X1_4
timestamp 1719641852
transform 1 0 3284 0 -1 1105
box -2 -3 50 103
use NOR2X1  NOR2X1_136
timestamp 1719641852
transform 1 0 3332 0 -1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_135
timestamp 1719641852
transform 1 0 3356 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_244
timestamp 1719641852
transform 1 0 3380 0 -1 1105
box -2 -3 34 103
use FILL  FILL_10_6_0
timestamp 1719641852
transform 1 0 3412 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_6_1
timestamp 1719641852
transform 1 0 3420 0 -1 1105
box -2 -3 10 103
use NOR2X1  NOR2X1_78
timestamp 1719641852
transform 1 0 3428 0 -1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_76
timestamp 1719641852
transform 1 0 3452 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_125
timestamp 1719641852
transform 1 0 3484 0 -1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_126
timestamp 1719641852
transform 1 0 3508 0 -1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_31
timestamp 1719641852
transform 1 0 3532 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_230
timestamp 1719641852
transform 1 0 3564 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_120
timestamp 1719641852
transform 1 0 3596 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_231
timestamp 1719641852
transform 1 0 3620 0 -1 1105
box -2 -3 34 103
use BUFX4  BUFX4_236
timestamp 1719641852
transform -1 0 3684 0 -1 1105
box -2 -3 34 103
use AND2X2  AND2X2_15
timestamp 1719641852
transform 1 0 3684 0 -1 1105
box -2 -3 34 103
use AND2X2  AND2X2_16
timestamp 1719641852
transform 1 0 3716 0 -1 1105
box -2 -3 34 103
use BUFX4  BUFX4_235
timestamp 1719641852
transform -1 0 3780 0 -1 1105
box -2 -3 34 103
use DFFSR  DFFSR_103
timestamp 1719641852
transform 1 0 4 0 1 1105
box -2 -3 178 103
use NOR2X1  NOR2X1_30
timestamp 1719641852
transform 1 0 180 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_163
timestamp 1719641852
transform -1 0 236 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_39
timestamp 1719641852
transform 1 0 236 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_165
timestamp 1719641852
transform -1 0 292 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_20
timestamp 1719641852
transform 1 0 292 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_161
timestamp 1719641852
transform -1 0 356 0 1 1105
box -2 -3 34 103
use FILL  FILL_11_0_0
timestamp 1719641852
transform 1 0 356 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_0_1
timestamp 1719641852
transform 1 0 364 0 1 1105
box -2 -3 10 103
use XOR2X1  XOR2X1_1
timestamp 1719641852
transform 1 0 372 0 1 1105
box -2 -3 58 103
use OAI21X1  OAI21X1_162
timestamp 1719641852
transform -1 0 460 0 1 1105
box -2 -3 34 103
use INVX2  INVX2_40
timestamp 1719641852
transform -1 0 476 0 1 1105
box -2 -3 18 103
use NAND2X1  NAND2X1_100
timestamp 1719641852
transform -1 0 500 0 1 1105
box -2 -3 26 103
use NAND3X1  NAND3X1_103
timestamp 1719641852
transform 1 0 500 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_32
timestamp 1719641852
transform -1 0 556 0 1 1105
box -2 -3 26 103
use BUFX4  BUFX4_104
timestamp 1719641852
transform -1 0 588 0 1 1105
box -2 -3 34 103
use INVX2  INVX2_29
timestamp 1719641852
transform 1 0 588 0 1 1105
box -2 -3 18 103
use DFFSR  DFFSR_101
timestamp 1719641852
transform -1 0 780 0 1 1105
box -2 -3 178 103
use INVX2  INVX2_3
timestamp 1719641852
transform 1 0 780 0 1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_38
timestamp 1719641852
transform 1 0 796 0 1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_21
timestamp 1719641852
transform 1 0 828 0 1 1105
box -2 -3 34 103
use FILL  FILL_11_1_0
timestamp 1719641852
transform -1 0 868 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_1_1
timestamp 1719641852
transform -1 0 876 0 1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_37
timestamp 1719641852
transform -1 0 908 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_19
timestamp 1719641852
transform -1 0 932 0 1 1105
box -2 -3 26 103
use BUFX4  BUFX4_17
timestamp 1719641852
transform -1 0 964 0 1 1105
box -2 -3 34 103
use BUFX4  BUFX4_14
timestamp 1719641852
transform -1 0 996 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_24
timestamp 1719641852
transform 1 0 996 0 1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_328
timestamp 1719641852
transform -1 0 1044 0 1 1105
box -2 -3 26 103
use OAI22X1  OAI22X1_25
timestamp 1719641852
transform 1 0 1044 0 1 1105
box -2 -3 42 103
use INVX1  INVX1_59
timestamp 1719641852
transform -1 0 1100 0 1 1105
box -2 -3 18 103
use OAI22X1  OAI22X1_36
timestamp 1719641852
transform 1 0 1100 0 1 1105
box -2 -3 42 103
use INVX1  INVX1_61
timestamp 1719641852
transform -1 0 1156 0 1 1105
box -2 -3 18 103
use DFFSR  DFFSR_163
timestamp 1719641852
transform -1 0 1332 0 1 1105
box -2 -3 178 103
use INVX2  INVX2_96
timestamp 1719641852
transform 1 0 1332 0 1 1105
box -2 -3 18 103
use NAND2X1  NAND2X1_313
timestamp 1719641852
transform 1 0 1348 0 1 1105
box -2 -3 26 103
use FILL  FILL_11_2_0
timestamp 1719641852
transform -1 0 1380 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_2_1
timestamp 1719641852
transform -1 0 1388 0 1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_707
timestamp 1719641852
transform -1 0 1420 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_236
timestamp 1719641852
transform -1 0 1444 0 1 1105
box -2 -3 26 103
use BUFX4  BUFX4_192
timestamp 1719641852
transform 1 0 1444 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_333
timestamp 1719641852
transform 1 0 1476 0 1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_260
timestamp 1719641852
transform -1 0 1532 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_21
timestamp 1719641852
transform 1 0 1532 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_769
timestamp 1719641852
transform 1 0 1556 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_258
timestamp 1719641852
transform -1 0 1620 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_303
timestamp 1719641852
transform 1 0 1620 0 1 1105
box -2 -3 26 103
use INVX8  INVX8_11
timestamp 1719641852
transform 1 0 1644 0 1 1105
box -2 -3 42 103
use CLKBUF1  CLKBUF1_39
timestamp 1719641852
transform 1 0 1684 0 1 1105
box -2 -3 74 103
use NOR2X1  NOR2X1_235
timestamp 1719641852
transform -1 0 1780 0 1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_214
timestamp 1719641852
transform -1 0 1812 0 1 1105
box -2 -3 34 103
use INVX8  INVX8_23
timestamp 1719641852
transform 1 0 1812 0 1 1105
box -2 -3 42 103
use INVX1  INVX1_53
timestamp 1719641852
transform -1 0 1868 0 1 1105
box -2 -3 18 103
use INVX2  INVX2_123
timestamp 1719641852
transform -1 0 1884 0 1 1105
box -2 -3 18 103
use FILL  FILL_11_3_0
timestamp 1719641852
transform -1 0 1892 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_3_1
timestamp 1719641852
transform -1 0 1900 0 1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_613
timestamp 1719641852
transform -1 0 1932 0 1 1105
box -2 -3 34 103
use DFFSR  DFFSR_159
timestamp 1719641852
transform -1 0 2108 0 1 1105
box -2 -3 178 103
use DFFSR  DFFSR_226
timestamp 1719641852
transform -1 0 2284 0 1 1105
box -2 -3 178 103
use OAI21X1  OAI21X1_522
timestamp 1719641852
transform -1 0 2316 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_181
timestamp 1719641852
transform 1 0 2316 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_519
timestamp 1719641852
transform -1 0 2380 0 1 1105
box -2 -3 34 103
use INVX4  INVX4_7
timestamp 1719641852
transform 1 0 2380 0 1 1105
box -2 -3 26 103
use FILL  FILL_11_4_0
timestamp 1719641852
transform 1 0 2404 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_4_1
timestamp 1719641852
transform 1 0 2412 0 1 1105
box -2 -3 10 103
use NOR2X1  NOR2X1_260
timestamp 1719641852
transform 1 0 2420 0 1 1105
box -2 -3 26 103
use INVX4  INVX4_8
timestamp 1719641852
transform -1 0 2468 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_520
timestamp 1719641852
transform 1 0 2468 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_383
timestamp 1719641852
transform -1 0 2532 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_125
timestamp 1719641852
transform 1 0 2532 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_126
timestamp 1719641852
transform 1 0 2564 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_218
timestamp 1719641852
transform 1 0 2596 0 1 1105
box -2 -3 26 103
use INVX1  INVX1_62
timestamp 1719641852
transform -1 0 2636 0 1 1105
box -2 -3 18 103
use DFFSR  DFFSR_221
timestamp 1719641852
transform -1 0 2812 0 1 1105
box -2 -3 178 103
use OAI21X1  OAI21X1_401
timestamp 1719641852
transform 1 0 2812 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_405
timestamp 1719641852
transform -1 0 2876 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_250
timestamp 1719641852
transform -1 0 2900 0 1 1105
box -2 -3 26 103
use FILL  FILL_11_5_0
timestamp 1719641852
transform -1 0 2908 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_5_1
timestamp 1719641852
transform -1 0 2916 0 1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_404
timestamp 1719641852
transform -1 0 2948 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_403
timestamp 1719641852
transform -1 0 2980 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_223
timestamp 1719641852
transform 1 0 2980 0 1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_133
timestamp 1719641852
transform 1 0 3004 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_402
timestamp 1719641852
transform 1 0 3036 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_206
timestamp 1719641852
transform 1 0 3068 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_389
timestamp 1719641852
transform 1 0 3092 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_387
timestamp 1719641852
transform 1 0 3124 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_202
timestamp 1719641852
transform -1 0 3180 0 1 1105
box -2 -3 26 103
use INVX1  INVX1_122
timestamp 1719641852
transform -1 0 3196 0 1 1105
box -2 -3 18 103
use MUX2X1  MUX2X1_2
timestamp 1719641852
transform -1 0 3244 0 1 1105
box -2 -3 50 103
use AOI21X1  AOI21X1_66
timestamp 1719641852
transform 1 0 3244 0 1 1105
box -2 -3 34 103
use AOI22X1  AOI22X1_45
timestamp 1719641852
transform -1 0 3316 0 1 1105
box -2 -3 42 103
use NAND2X1  NAND2X1_167
timestamp 1719641852
transform -1 0 3340 0 1 1105
box -2 -3 26 103
use MUX2X1  MUX2X1_1
timestamp 1719641852
transform 1 0 3340 0 1 1105
box -2 -3 50 103
use NOR2X1  NOR2X1_76
timestamp 1719641852
transform 1 0 3388 0 1 1105
box -2 -3 26 103
use FILL  FILL_11_6_0
timestamp 1719641852
transform 1 0 3412 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_6_1
timestamp 1719641852
transform 1 0 3420 0 1 1105
box -2 -3 10 103
use NOR2X1  NOR2X1_75
timestamp 1719641852
transform 1 0 3428 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_208
timestamp 1719641852
transform 1 0 3452 0 1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_203
timestamp 1719641852
transform -1 0 3516 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_77
timestamp 1719641852
transform 1 0 3516 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_209
timestamp 1719641852
transform 1 0 3540 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_119
timestamp 1719641852
transform 1 0 3572 0 1 1105
box -2 -3 26 103
use NAND3X1  NAND3X1_113
timestamp 1719641852
transform -1 0 3628 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_118
timestamp 1719641852
transform 1 0 3628 0 1 1105
box -2 -3 26 103
use BUFX4  BUFX4_238
timestamp 1719641852
transform -1 0 3684 0 1 1105
box -2 -3 34 103
use BUFX4  BUFX4_195
timestamp 1719641852
transform 1 0 3684 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_232
timestamp 1719641852
transform 1 0 3716 0 1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_133
timestamp 1719641852
transform -1 0 3780 0 1 1105
box -2 -3 34 103
use BUFX4  BUFX4_88
timestamp 1719641852
transform -1 0 36 0 -1 1305
box -2 -3 34 103
use CLKBUF1  CLKBUF1_63
timestamp 1719641852
transform 1 0 36 0 -1 1305
box -2 -3 74 103
use CLKBUF1  CLKBUF1_21
timestamp 1719641852
transform -1 0 180 0 -1 1305
box -2 -3 74 103
use INVX1  INVX1_70
timestamp 1719641852
transform 1 0 180 0 -1 1305
box -2 -3 18 103
use NAND2X1  NAND2X1_89
timestamp 1719641852
transform 1 0 196 0 -1 1305
box -2 -3 26 103
use AND2X2  AND2X2_6
timestamp 1719641852
transform 1 0 220 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_91
timestamp 1719641852
transform -1 0 276 0 -1 1305
box -2 -3 26 103
use FILL  FILL_12_0_0
timestamp 1719641852
transform -1 0 284 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_0_1
timestamp 1719641852
transform -1 0 292 0 -1 1305
box -2 -3 10 103
use DFFSR  DFFSR_99
timestamp 1719641852
transform -1 0 468 0 -1 1305
box -2 -3 178 103
use INVX1  INVX1_66
timestamp 1719641852
transform 1 0 468 0 -1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_159
timestamp 1719641852
transform 1 0 484 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_85
timestamp 1719641852
transform -1 0 540 0 -1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_83
timestamp 1719641852
transform -1 0 564 0 -1 1305
box -2 -3 26 103
use OR2X2  OR2X2_3
timestamp 1719641852
transform -1 0 596 0 -1 1305
box -2 -3 34 103
use DFFSR  DFFSR_62
timestamp 1719641852
transform -1 0 772 0 -1 1305
box -2 -3 178 103
use INVX2  INVX2_30
timestamp 1719641852
transform 1 0 772 0 -1 1305
box -2 -3 18 103
use FILL  FILL_12_1_0
timestamp 1719641852
transform 1 0 788 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_1_1
timestamp 1719641852
transform 1 0 796 0 -1 1305
box -2 -3 10 103
use DFFSR  DFFSR_56
timestamp 1719641852
transform 1 0 804 0 -1 1305
box -2 -3 178 103
use NOR2X1  NOR2X1_1
timestamp 1719641852
transform 1 0 980 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_108
timestamp 1719641852
transform -1 0 1036 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_14
timestamp 1719641852
transform -1 0 1060 0 -1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_53
timestamp 1719641852
transform -1 0 1084 0 -1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_11
timestamp 1719641852
transform -1 0 1116 0 -1 1305
box -2 -3 34 103
use OAI22X1  OAI22X1_37
timestamp 1719641852
transform 1 0 1116 0 -1 1305
box -2 -3 42 103
use AOI21X1  AOI21X1_17
timestamp 1719641852
transform -1 0 1188 0 -1 1305
box -2 -3 34 103
use DFFSR  DFFSR_161
timestamp 1719641852
transform 1 0 1188 0 -1 1305
box -2 -3 178 103
use FILL  FILL_12_2_0
timestamp 1719641852
transform -1 0 1372 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_2_1
timestamp 1719641852
transform -1 0 1380 0 -1 1305
box -2 -3 10 103
use INVX1  INVX1_57
timestamp 1719641852
transform -1 0 1396 0 -1 1305
box -2 -3 18 103
use INVX2  INVX2_154
timestamp 1719641852
transform 1 0 1396 0 -1 1305
box -2 -3 18 103
use NOR2X1  NOR2X1_284
timestamp 1719641852
transform 1 0 1412 0 -1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_218
timestamp 1719641852
transform -1 0 1468 0 -1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_217
timestamp 1719641852
transform -1 0 1500 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_615
timestamp 1719641852
transform -1 0 1532 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_155
timestamp 1719641852
transform 1 0 1532 0 -1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_614
timestamp 1719641852
transform 1 0 1548 0 -1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_216
timestamp 1719641852
transform -1 0 1612 0 -1 1305
box -2 -3 34 103
use BUFX4  BUFX4_96
timestamp 1719641852
transform -1 0 1644 0 -1 1305
box -2 -3 34 103
use CLKBUF1  CLKBUF1_67
timestamp 1719641852
transform -1 0 1716 0 -1 1305
box -2 -3 74 103
use INVX1  INVX1_146
timestamp 1719641852
transform -1 0 1732 0 -1 1305
box -2 -3 18 103
use NAND2X1  NAND2X1_311
timestamp 1719641852
transform -1 0 1756 0 -1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_276
timestamp 1719641852
transform -1 0 1780 0 -1 1305
box -2 -3 26 103
use BUFX4  BUFX4_64
timestamp 1719641852
transform -1 0 1812 0 -1 1305
box -2 -3 34 103
use FILL  FILL_12_3_0
timestamp 1719641852
transform -1 0 1820 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_3_1
timestamp 1719641852
transform -1 0 1828 0 -1 1305
box -2 -3 10 103
use DFFSR  DFFSR_192
timestamp 1719641852
transform -1 0 2004 0 -1 1305
box -2 -3 178 103
use NOR2X1  NOR2X1_302
timestamp 1719641852
transform -1 0 2028 0 -1 1305
box -2 -3 26 103
use BUFX4  BUFX4_30
timestamp 1719641852
transform -1 0 2060 0 -1 1305
box -2 -3 34 103
use DFFSR  DFFSR_188
timestamp 1719641852
transform -1 0 2236 0 -1 1305
box -2 -3 178 103
use AOI21X1  AOI21X1_219
timestamp 1719641852
transform 1 0 2236 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_616
timestamp 1719641852
transform -1 0 2300 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_518
timestamp 1719641852
transform -1 0 2332 0 -1 1305
box -2 -3 34 103
use INVX2  INVX2_98
timestamp 1719641852
transform 1 0 2332 0 -1 1305
box -2 -3 18 103
use AOI21X1  AOI21X1_174
timestamp 1719641852
transform -1 0 2380 0 -1 1305
box -2 -3 34 103
use FILL  FILL_12_4_0
timestamp 1719641852
transform -1 0 2388 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_4_1
timestamp 1719641852
transform -1 0 2396 0 -1 1305
box -2 -3 10 103
use OAI21X1  OAI21X1_498
timestamp 1719641852
transform -1 0 2428 0 -1 1305
box -2 -3 34 103
use BUFX4  BUFX4_119
timestamp 1719641852
transform 1 0 2428 0 -1 1305
box -2 -3 34 103
use BUFX4  BUFX4_167
timestamp 1719641852
transform 1 0 2460 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_256
timestamp 1719641852
transform 1 0 2492 0 -1 1305
box -2 -3 26 103
use BUFX4  BUFX4_129
timestamp 1719641852
transform 1 0 2516 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_257
timestamp 1719641852
transform 1 0 2548 0 -1 1305
box -2 -3 26 103
use BUFX4  BUFX4_99
timestamp 1719641852
transform 1 0 2572 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_575
timestamp 1719641852
transform 1 0 2604 0 -1 1305
box -2 -3 34 103
use DFFSR  DFFSR_220
timestamp 1719641852
transform -1 0 2812 0 -1 1305
box -2 -3 178 103
use INVX2  INVX2_99
timestamp 1719641852
transform 1 0 2812 0 -1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_443
timestamp 1719641852
transform 1 0 2828 0 -1 1305
box -2 -3 34 103
use BUFX4  BUFX4_148
timestamp 1719641852
transform -1 0 2892 0 -1 1305
box -2 -3 34 103
use FILL  FILL_12_5_0
timestamp 1719641852
transform -1 0 2900 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_5_1
timestamp 1719641852
transform -1 0 2908 0 -1 1305
box -2 -3 10 103
use BUFX4  BUFX4_243
timestamp 1719641852
transform -1 0 2940 0 -1 1305
box -2 -3 34 103
use INVX2  INVX2_140
timestamp 1719641852
transform 1 0 2940 0 -1 1305
box -2 -3 18 103
use NOR2X1  NOR2X1_201
timestamp 1719641852
transform 1 0 2956 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_438
timestamp 1719641852
transform 1 0 2980 0 -1 1305
box -2 -3 34 103
use INVX8  INVX8_16
timestamp 1719641852
transform 1 0 3012 0 -1 1305
box -2 -3 42 103
use OAI21X1  OAI21X1_386
timestamp 1719641852
transform -1 0 3084 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_124
timestamp 1719641852
transform -1 0 3100 0 -1 1305
box -2 -3 18 103
use BUFX4  BUFX4_54
timestamp 1719641852
transform 1 0 3100 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_392
timestamp 1719641852
transform 1 0 3132 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_393
timestamp 1719641852
transform 1 0 3164 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_205
timestamp 1719641852
transform -1 0 3220 0 -1 1305
box -2 -3 26 103
use INVX1  INVX1_123
timestamp 1719641852
transform -1 0 3236 0 -1 1305
box -2 -3 18 103
use INVX8  INVX8_17
timestamp 1719641852
transform 1 0 3236 0 -1 1305
box -2 -3 42 103
use AOI21X1  AOI21X1_63
timestamp 1719641852
transform 1 0 3276 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_169
timestamp 1719641852
transform -1 0 3332 0 -1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_82
timestamp 1719641852
transform 1 0 3332 0 -1 1305
box -2 -3 34 103
use AOI22X1  AOI22X1_53
timestamp 1719641852
transform -1 0 3404 0 -1 1305
box -2 -3 42 103
use NAND2X1  NAND2X1_183
timestamp 1719641852
transform -1 0 3428 0 -1 1305
box -2 -3 26 103
use FILL  FILL_12_6_0
timestamp 1719641852
transform -1 0 3436 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_6_1
timestamp 1719641852
transform -1 0 3444 0 -1 1305
box -2 -3 10 103
use AOI22X1  AOI22X1_49
timestamp 1719641852
transform -1 0 3484 0 -1 1305
box -2 -3 42 103
use NAND2X1  NAND2X1_184
timestamp 1719641852
transform -1 0 3508 0 -1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_123
timestamp 1719641852
transform 1 0 3508 0 -1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_30
timestamp 1719641852
transform 1 0 3532 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_124
timestamp 1719641852
transform 1 0 3564 0 -1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_157
timestamp 1719641852
transform 1 0 3588 0 -1 1305
box -2 -3 26 103
use NAND3X1  NAND3X1_115
timestamp 1719641852
transform -1 0 3644 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_160
timestamp 1719641852
transform -1 0 3668 0 -1 1305
box -2 -3 26 103
use AOI22X1  AOI22X1_39
timestamp 1719641852
transform -1 0 3708 0 -1 1305
box -2 -3 42 103
use AOI21X1  AOI21X1_56
timestamp 1719641852
transform -1 0 3740 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_156
timestamp 1719641852
transform -1 0 3764 0 -1 1305
box -2 -3 26 103
use FILL  FILL_13_1
timestamp 1719641852
transform -1 0 3772 0 -1 1305
box -2 -3 10 103
use FILL  FILL_13_2
timestamp 1719641852
transform -1 0 3780 0 -1 1305
box -2 -3 10 103
use INVX8  INVX8_8
timestamp 1719641852
transform -1 0 44 0 1 1305
box -2 -3 42 103
use BUFX2  BUFX2_46
timestamp 1719641852
transform -1 0 68 0 1 1305
box -2 -3 26 103
use DFFSR  DFFSR_75
timestamp 1719641852
transform -1 0 244 0 1 1305
box -2 -3 178 103
use OAI21X1  OAI21X1_164
timestamp 1719641852
transform 1 0 244 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_92
timestamp 1719641852
transform -1 0 300 0 1 1305
box -2 -3 26 103
use FILL  FILL_13_0_0
timestamp 1719641852
transform 1 0 300 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_0_1
timestamp 1719641852
transform 1 0 308 0 1 1305
box -2 -3 10 103
use DFFSR  DFFSR_58
timestamp 1719641852
transform 1 0 316 0 1 1305
box -2 -3 178 103
use INVX1  INVX1_69
timestamp 1719641852
transform -1 0 508 0 1 1305
box -2 -3 18 103
use NOR2X1  NOR2X1_34
timestamp 1719641852
transform 1 0 508 0 1 1305
box -2 -3 26 103
use NAND3X1  NAND3X1_104
timestamp 1719641852
transform 1 0 532 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_33
timestamp 1719641852
transform 1 0 564 0 1 1305
box -2 -3 26 103
use INVX8  INVX8_7
timestamp 1719641852
transform 1 0 588 0 1 1305
box -2 -3 42 103
use INVX8  INVX8_24
timestamp 1719641852
transform 1 0 628 0 1 1305
box -2 -3 42 103
use OAI21X1  OAI21X1_107
timestamp 1719641852
transform 1 0 668 0 1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_57
timestamp 1719641852
transform 1 0 700 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_106
timestamp 1719641852
transform -1 0 764 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_109
timestamp 1719641852
transform 1 0 764 0 1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_58
timestamp 1719641852
transform -1 0 828 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_97
timestamp 1719641852
transform 1 0 828 0 1 1305
box -2 -3 34 103
use FILL  FILL_13_1_0
timestamp 1719641852
transform -1 0 868 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_1_1
timestamp 1719641852
transform -1 0 876 0 1 1305
box -2 -3 10 103
use AND2X2  AND2X2_1
timestamp 1719641852
transform -1 0 908 0 1 1305
box -2 -3 34 103
use INVX2  INVX2_24
timestamp 1719641852
transform -1 0 924 0 1 1305
box -2 -3 18 103
use NAND2X1  NAND2X1_231
timestamp 1719641852
transform 1 0 924 0 1 1305
box -2 -3 26 103
use OAI22X1  OAI22X1_26
timestamp 1719641852
transform 1 0 948 0 1 1305
box -2 -3 42 103
use INVX1  INVX1_51
timestamp 1719641852
transform -1 0 1004 0 1 1305
box -2 -3 18 103
use DFFSR  DFFSR_129
timestamp 1719641852
transform 1 0 1004 0 1 1305
box -2 -3 178 103
use DFFSR  DFFSR_193
timestamp 1719641852
transform 1 0 1180 0 1 1305
box -2 -3 178 103
use INVX1  INVX1_58
timestamp 1719641852
transform -1 0 1372 0 1 1305
box -2 -3 18 103
use FILL  FILL_13_2_0
timestamp 1719641852
transform 1 0 1372 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_2_1
timestamp 1719641852
transform 1 0 1380 0 1 1305
box -2 -3 10 103
use NAND2X1  NAND2X1_307
timestamp 1719641852
transform 1 0 1388 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_698
timestamp 1719641852
transform -1 0 1444 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_696
timestamp 1719641852
transform -1 0 1476 0 1 1305
box -2 -3 34 103
use INVX2  INVX2_156
timestamp 1719641852
transform -1 0 1492 0 1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_697
timestamp 1719641852
transform -1 0 1524 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_317
timestamp 1719641852
transform -1 0 1548 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_706
timestamp 1719641852
transform -1 0 1580 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_312
timestamp 1719641852
transform 1 0 1580 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_705
timestamp 1719641852
transform -1 0 1636 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_704
timestamp 1719641852
transform 1 0 1636 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_703
timestamp 1719641852
transform -1 0 1700 0 1 1305
box -2 -3 34 103
use OAI22X1  OAI22X1_28
timestamp 1719641852
transform 1 0 1700 0 1 1305
box -2 -3 42 103
use AOI21X1  AOI21X1_227
timestamp 1719641852
transform -1 0 1772 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_628
timestamp 1719641852
transform -1 0 1804 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_626
timestamp 1719641852
transform -1 0 1836 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_625
timestamp 1719641852
transform -1 0 1868 0 1 1305
box -2 -3 34 103
use INVX1  INVX1_52
timestamp 1719641852
transform -1 0 1884 0 1 1305
box -2 -3 18 103
use FILL  FILL_13_3_0
timestamp 1719641852
transform -1 0 1892 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_3_1
timestamp 1719641852
transform -1 0 1900 0 1 1305
box -2 -3 10 103
use DFFSR  DFFSR_160
timestamp 1719641852
transform -1 0 2076 0 1 1305
box -2 -3 178 103
use NAND2X1  NAND2X1_272
timestamp 1719641852
transform 1 0 2076 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_619
timestamp 1719641852
transform -1 0 2132 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_618
timestamp 1719641852
transform -1 0 2164 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_617
timestamp 1719641852
transform -1 0 2196 0 1 1305
box -2 -3 34 103
use BUFX4  BUFX4_120
timestamp 1719641852
transform -1 0 2228 0 1 1305
box -2 -3 34 103
use INVX1  INVX1_54
timestamp 1719641852
transform -1 0 2244 0 1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_497
timestamp 1719641852
transform 1 0 2244 0 1 1305
box -2 -3 34 103
use INVX2  INVX2_155
timestamp 1719641852
transform 1 0 2276 0 1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_501
timestamp 1719641852
transform -1 0 2324 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_500
timestamp 1719641852
transform -1 0 2356 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_499
timestamp 1719641852
transform -1 0 2388 0 1 1305
box -2 -3 34 103
use FILL  FILL_13_4_0
timestamp 1719641852
transform 1 0 2388 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_4_1
timestamp 1719641852
transform 1 0 2396 0 1 1305
box -2 -3 10 103
use OAI21X1  OAI21X1_502
timestamp 1719641852
transform 1 0 2404 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_506
timestamp 1719641852
transform -1 0 2468 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_505
timestamp 1719641852
transform -1 0 2500 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_504
timestamp 1719641852
transform -1 0 2532 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_503
timestamp 1719641852
transform -1 0 2564 0 1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_175
timestamp 1719641852
transform -1 0 2596 0 1 1305
box -2 -3 34 103
use DFFSR  DFFSR_235
timestamp 1719641852
transform -1 0 2772 0 1 1305
box -2 -3 178 103
use OAI21X1  OAI21X1_410
timestamp 1719641852
transform -1 0 2804 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_408
timestamp 1719641852
transform -1 0 2836 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_409
timestamp 1719641852
transform -1 0 2868 0 1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_134
timestamp 1719641852
transform 1 0 2868 0 1 1305
box -2 -3 34 103
use FILL  FILL_13_5_0
timestamp 1719641852
transform -1 0 2908 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_5_1
timestamp 1719641852
transform -1 0 2916 0 1 1305
box -2 -3 10 103
use OAI21X1  OAI21X1_407
timestamp 1719641852
transform -1 0 2948 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_224
timestamp 1719641852
transform 1 0 2948 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_391
timestamp 1719641852
transform -1 0 3004 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_390
timestamp 1719641852
transform -1 0 3036 0 1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_128
timestamp 1719641852
transform -1 0 3068 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_220
timestamp 1719641852
transform -1 0 3092 0 1 1305
box -2 -3 26 103
use INVX2  INVX2_164
timestamp 1719641852
transform -1 0 3108 0 1 1305
box -2 -3 18 103
use INVX2  INVX2_84
timestamp 1719641852
transform 1 0 3108 0 1 1305
box -2 -3 18 103
use NAND2X1  NAND2X1_211
timestamp 1719641852
transform 1 0 3124 0 1 1305
box -2 -3 26 103
use BUFX4  BUFX4_67
timestamp 1719641852
transform -1 0 3180 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_203
timestamp 1719641852
transform -1 0 3204 0 1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_64
timestamp 1719641852
transform 1 0 3204 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_166
timestamp 1719641852
transform 1 0 3236 0 1 1305
box -2 -3 26 103
use AOI22X1  AOI22X1_44
timestamp 1719641852
transform -1 0 3300 0 1 1305
box -2 -3 42 103
use NAND2X1  NAND2X1_165
timestamp 1719641852
transform -1 0 3324 0 1 1305
box -2 -3 26 103
use INVX2  INVX2_86
timestamp 1719641852
transform -1 0 3340 0 1 1305
box -2 -3 18 103
use AOI21X1  AOI21X1_81
timestamp 1719641852
transform 1 0 3340 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_176
timestamp 1719641852
transform 1 0 3372 0 1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_75
timestamp 1719641852
transform 1 0 3396 0 1 1305
box -2 -3 34 103
use FILL  FILL_13_6_0
timestamp 1719641852
transform 1 0 3428 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_6_1
timestamp 1719641852
transform 1 0 3436 0 1 1305
box -2 -3 10 103
use NAND3X1  NAND3X1_202
timestamp 1719641852
transform 1 0 3444 0 1 1305
box -2 -3 34 103
use BUFX4  BUFX4_153
timestamp 1719641852
transform -1 0 3508 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_164
timestamp 1719641852
transform 1 0 3508 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_252
timestamp 1719641852
transform 1 0 3532 0 1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_57
timestamp 1719641852
transform 1 0 3564 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_165
timestamp 1719641852
transform 1 0 3596 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_260
timestamp 1719641852
transform 1 0 3620 0 1 1305
box -2 -3 34 103
use BUFX4  BUFX4_158
timestamp 1719641852
transform 1 0 3652 0 1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_161
timestamp 1719641852
transform -1 0 3716 0 1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_162
timestamp 1719641852
transform -1 0 3748 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_259
timestamp 1719641852
transform 1 0 3748 0 1 1305
box -2 -3 34 103
use DFFSR  DFFSR_102
timestamp 1719641852
transform 1 0 4 0 -1 1505
box -2 -3 178 103
use DFFSR  DFFSR_97
timestamp 1719641852
transform 1 0 180 0 -1 1505
box -2 -3 178 103
use FILL  FILL_14_0_0
timestamp 1719641852
transform -1 0 364 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_0_1
timestamp 1719641852
transform -1 0 372 0 -1 1505
box -2 -3 10 103
use INVX1  INVX1_67
timestamp 1719641852
transform -1 0 388 0 -1 1505
box -2 -3 18 103
use OAI22X1  OAI22X1_40
timestamp 1719641852
transform -1 0 428 0 -1 1505
box -2 -3 42 103
use OR2X2  OR2X2_1
timestamp 1719641852
transform -1 0 460 0 -1 1505
box -2 -3 34 103
use OAI22X1  OAI22X1_41
timestamp 1719641852
transform -1 0 500 0 -1 1505
box -2 -3 42 103
use INVX2  INVX2_26
timestamp 1719641852
transform 1 0 500 0 -1 1505
box -2 -3 18 103
use INVX1  INVX1_68
timestamp 1719641852
transform 1 0 516 0 -1 1505
box -2 -3 18 103
use INVX2  INVX2_25
timestamp 1719641852
transform 1 0 532 0 -1 1505
box -2 -3 18 103
use DFFSR  DFFSR_98
timestamp 1719641852
transform 1 0 548 0 -1 1505
box -2 -3 178 103
use NAND2X1  NAND2X1_23
timestamp 1719641852
transform -1 0 748 0 -1 1505
box -2 -3 26 103
use BUFX4  BUFX4_5
timestamp 1719641852
transform 1 0 748 0 -1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_52
timestamp 1719641852
transform -1 0 812 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_96
timestamp 1719641852
transform -1 0 844 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_18
timestamp 1719641852
transform -1 0 868 0 -1 1505
box -2 -3 26 103
use FILL  FILL_14_1_0
timestamp 1719641852
transform -1 0 876 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_1_1
timestamp 1719641852
transform -1 0 884 0 -1 1505
box -2 -3 10 103
use BUFX4  BUFX4_6
timestamp 1719641852
transform -1 0 916 0 -1 1505
box -2 -3 34 103
use BUFX4  BUFX4_12
timestamp 1719641852
transform 1 0 916 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_237
timestamp 1719641852
transform -1 0 972 0 -1 1505
box -2 -3 26 103
use OAI22X1  OAI22X1_24
timestamp 1719641852
transform 1 0 972 0 -1 1505
box -2 -3 42 103
use NAND2X1  NAND2X1_20
timestamp 1719641852
transform 1 0 1012 0 -1 1505
box -2 -3 26 103
use INVX1  INVX1_49
timestamp 1719641852
transform -1 0 1052 0 -1 1505
box -2 -3 18 103
use OAI22X1  OAI22X1_34
timestamp 1719641852
transform -1 0 1092 0 -1 1505
box -2 -3 42 103
use AOI21X1  AOI21X1_14
timestamp 1719641852
transform -1 0 1124 0 -1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_12
timestamp 1719641852
transform 1 0 1124 0 -1 1505
box -2 -3 34 103
use OAI22X1  OAI22X1_29
timestamp 1719641852
transform 1 0 1156 0 -1 1505
box -2 -3 42 103
use BUFX4  BUFX4_190
timestamp 1719641852
transform -1 0 1228 0 -1 1505
box -2 -3 34 103
use CLKBUF1  CLKBUF1_1
timestamp 1719641852
transform 1 0 1228 0 -1 1505
box -2 -3 74 103
use OAI22X1  OAI22X1_33
timestamp 1719641852
transform 1 0 1300 0 -1 1505
box -2 -3 42 103
use FILL  FILL_14_2_0
timestamp 1719641852
transform -1 0 1348 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_2_1
timestamp 1719641852
transform -1 0 1356 0 -1 1505
box -2 -3 10 103
use DFFSR  DFFSR_125
timestamp 1719641852
transform -1 0 1532 0 -1 1505
box -2 -3 178 103
use INVX2  INVX2_138
timestamp 1719641852
transform 1 0 1532 0 -1 1505
box -2 -3 18 103
use DFFSR  DFFSR_157
timestamp 1719641852
transform -1 0 1724 0 -1 1505
box -2 -3 178 103
use INVX2  INVX2_136
timestamp 1719641852
transform 1 0 1724 0 -1 1505
box -2 -3 18 103
use INVX2  INVX2_97
timestamp 1719641852
transform 1 0 1740 0 -1 1505
box -2 -3 18 103
use NAND2X1  NAND2X1_275
timestamp 1719641852
transform 1 0 1756 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_627
timestamp 1719641852
transform -1 0 1812 0 -1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_226
timestamp 1719641852
transform 1 0 1812 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_624
timestamp 1719641852
transform -1 0 1876 0 -1 1505
box -2 -3 34 103
use FILL  FILL_14_3_0
timestamp 1719641852
transform -1 0 1884 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_3_1
timestamp 1719641852
transform -1 0 1892 0 -1 1505
box -2 -3 10 103
use OAI21X1  OAI21X1_629
timestamp 1719641852
transform -1 0 1924 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_287
timestamp 1719641852
transform -1 0 1948 0 -1 1505
box -2 -3 26 103
use DFFSR  DFFSR_217
timestamp 1719641852
transform -1 0 2124 0 -1 1505
box -2 -3 178 103
use INVX2  INVX2_85
timestamp 1719641852
transform 1 0 2124 0 -1 1505
box -2 -3 18 103
use DFFSR  DFFSR_189
timestamp 1719641852
transform -1 0 2316 0 -1 1505
box -2 -3 178 103
use OAI21X1  OAI21X1_513
timestamp 1719641852
transform 1 0 2316 0 -1 1505
box -2 -3 34 103
use INVX2  INVX2_142
timestamp 1719641852
transform 1 0 2348 0 -1 1505
box -2 -3 18 103
use OAI21X1  OAI21X1_517
timestamp 1719641852
transform -1 0 2396 0 -1 1505
box -2 -3 34 103
use FILL  FILL_14_4_0
timestamp 1719641852
transform -1 0 2404 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_4_1
timestamp 1719641852
transform -1 0 2412 0 -1 1505
box -2 -3 10 103
use OAI21X1  OAI21X1_516
timestamp 1719641852
transform -1 0 2444 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_515
timestamp 1719641852
transform -1 0 2476 0 -1 1505
box -2 -3 34 103
use BUFX4  BUFX4_166
timestamp 1719641852
transform 1 0 2476 0 -1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_180
timestamp 1719641852
transform 1 0 2508 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_514
timestamp 1719641852
transform -1 0 2572 0 -1 1505
box -2 -3 34 103
use INVX4  INVX4_9
timestamp 1719641852
transform -1 0 2596 0 -1 1505
box -2 -3 26 103
use INVX4  INVX4_10
timestamp 1719641852
transform 1 0 2596 0 -1 1505
box -2 -3 26 103
use AND2X2  AND2X2_24
timestamp 1719641852
transform -1 0 2652 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_746
timestamp 1719641852
transform -1 0 2684 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_750
timestamp 1719641852
transform -1 0 2716 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_749
timestamp 1719641852
transform -1 0 2748 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_406
timestamp 1719641852
transform 1 0 2748 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_416
timestamp 1719641852
transform -1 0 2812 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_420
timestamp 1719641852
transform -1 0 2844 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_419
timestamp 1719641852
transform 1 0 2844 0 -1 1505
box -2 -3 34 103
use BUFX4  BUFX4_221
timestamp 1719641852
transform -1 0 2908 0 -1 1505
box -2 -3 34 103
use FILL  FILL_14_5_0
timestamp 1719641852
transform 1 0 2908 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_5_1
timestamp 1719641852
transform 1 0 2916 0 -1 1505
box -2 -3 10 103
use BUFX4  BUFX4_220
timestamp 1719641852
transform 1 0 2924 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_239
timestamp 1719641852
transform 1 0 2956 0 -1 1505
box -2 -3 26 103
use BUFX4  BUFX4_149
timestamp 1719641852
transform 1 0 2980 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_209
timestamp 1719641852
transform -1 0 3036 0 -1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_193
timestamp 1719641852
transform -1 0 3060 0 -1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_197
timestamp 1719641852
transform 1 0 3060 0 -1 1505
box -2 -3 26 103
use BUFX4  BUFX4_51
timestamp 1719641852
transform 1 0 3084 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_196
timestamp 1719641852
transform -1 0 3140 0 -1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_182
timestamp 1719641852
transform -1 0 3164 0 -1 1505
box -2 -3 26 103
use INVX1  INVX1_126
timestamp 1719641852
transform -1 0 3180 0 -1 1505
box -2 -3 18 103
use INVX1  INVX1_125
timestamp 1719641852
transform -1 0 3196 0 -1 1505
box -2 -3 18 103
use AOI21X1  AOI21X1_102
timestamp 1719641852
transform 1 0 3196 0 -1 1505
box -2 -3 34 103
use INVX1  INVX1_121
timestamp 1719641852
transform 1 0 3228 0 -1 1505
box -2 -3 18 103
use NOR2X1  NOR2X1_200
timestamp 1719641852
transform -1 0 3268 0 -1 1505
box -2 -3 26 103
use NOR3X1  NOR3X1_3
timestamp 1719641852
transform 1 0 3268 0 -1 1505
box -2 -3 66 103
use BUFX4  BUFX4_155
timestamp 1719641852
transform -1 0 3364 0 -1 1505
box -2 -3 34 103
use BUFX4  BUFX4_173
timestamp 1719641852
transform 1 0 3364 0 -1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_85
timestamp 1719641852
transform -1 0 3428 0 -1 1505
box -2 -3 34 103
use FILL  FILL_14_6_0
timestamp 1719641852
transform 1 0 3428 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_6_1
timestamp 1719641852
transform 1 0 3436 0 -1 1505
box -2 -3 10 103
use OAI21X1  OAI21X1_299
timestamp 1719641852
transform 1 0 3444 0 -1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_73
timestamp 1719641852
transform -1 0 3508 0 -1 1505
box -2 -3 34 103
use BUFX4  BUFX4_175
timestamp 1719641852
transform -1 0 3540 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_102
timestamp 1719641852
transform 1 0 3540 0 -1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_101
timestamp 1719641852
transform 1 0 3564 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_221
timestamp 1719641852
transform 1 0 3588 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_103
timestamp 1719641852
transform 1 0 3620 0 -1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_104
timestamp 1719641852
transform 1 0 3644 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_222
timestamp 1719641852
transform 1 0 3668 0 -1 1505
box -2 -3 34 103
use BUFX4  BUFX4_177
timestamp 1719641852
transform 1 0 3700 0 -1 1505
box -2 -3 34 103
use BUFX4  BUFX4_188
timestamp 1719641852
transform -1 0 3764 0 -1 1505
box -2 -3 34 103
use FILL  FILL_15_1
timestamp 1719641852
transform -1 0 3772 0 -1 1505
box -2 -3 10 103
use FILL  FILL_15_2
timestamp 1719641852
transform -1 0 3780 0 -1 1505
box -2 -3 10 103
use BUFX2  BUFX2_49
timestamp 1719641852
transform -1 0 28 0 1 1505
box -2 -3 26 103
use BUFX2  BUFX2_2
timestamp 1719641852
transform -1 0 52 0 1 1505
box -2 -3 26 103
use CLKBUF1  CLKBUF1_25
timestamp 1719641852
transform -1 0 124 0 1 1505
box -2 -3 74 103
use DFFSR  DFFSR_59
timestamp 1719641852
transform 1 0 124 0 1 1505
box -2 -3 178 103
use DFFSR  DFFSR_78
timestamp 1719641852
transform -1 0 180 0 -1 1705
box -2 -3 178 103
use DFFSR  DFFSR_57
timestamp 1719641852
transform 1 0 180 0 -1 1705
box -2 -3 178 103
use NAND2X1  NAND2X1_90
timestamp 1719641852
transform -1 0 324 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_87
timestamp 1719641852
transform -1 0 348 0 1 1505
box -2 -3 26 103
use FILL  FILL_15_0_0
timestamp 1719641852
transform 1 0 348 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_0_1
timestamp 1719641852
transform 1 0 356 0 1 1505
box -2 -3 10 103
use NAND2X1  NAND2X1_88
timestamp 1719641852
transform 1 0 364 0 1 1505
box -2 -3 26 103
use FILL  FILL_16_0_0
timestamp 1719641852
transform -1 0 364 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_0_1
timestamp 1719641852
transform -1 0 372 0 -1 1705
box -2 -3 10 103
use NAND2X1  NAND2X1_82
timestamp 1719641852
transform -1 0 412 0 1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_19
timestamp 1719641852
transform -1 0 444 0 1 1505
box -2 -3 34 103
use INVX2  INVX2_27
timestamp 1719641852
transform 1 0 444 0 1 1505
box -2 -3 18 103
use OAI21X1  OAI21X1_103
timestamp 1719641852
transform 1 0 460 0 1 1505
box -2 -3 34 103
use BUFX4  BUFX4_8
timestamp 1719641852
transform 1 0 492 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_101
timestamp 1719641852
transform 1 0 524 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_37
timestamp 1719641852
transform -1 0 396 0 -1 1705
box -2 -3 26 103
use DFFSR  DFFSR_60
timestamp 1719641852
transform -1 0 572 0 -1 1705
box -2 -3 178 103
use NAND2X1  NAND2X1_22
timestamp 1719641852
transform -1 0 596 0 -1 1705
box -2 -3 26 103
use NAND3X1  NAND3X1_55
timestamp 1719641852
transform -1 0 588 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_99
timestamp 1719641852
transform 1 0 596 0 -1 1705
box -2 -3 34 103
use BUFX4  BUFX4_7
timestamp 1719641852
transform 1 0 620 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_102
timestamp 1719641852
transform -1 0 620 0 1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_53
timestamp 1719641852
transform 1 0 628 0 -1 1705
box -2 -3 34 103
use BUFX4  BUFX4_108
timestamp 1719641852
transform 1 0 652 0 1 1505
box -2 -3 34 103
use BUFX4  BUFX4_105
timestamp 1719641852
transform -1 0 716 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_21
timestamp 1719641852
transform 1 0 660 0 -1 1705
box -2 -3 26 103
use NAND3X1  NAND3X1_54
timestamp 1719641852
transform 1 0 684 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_98
timestamp 1719641852
transform 1 0 716 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_100
timestamp 1719641852
transform 1 0 716 0 1 1505
box -2 -3 34 103
use OAI22X1  OAI22X1_27
timestamp 1719641852
transform -1 0 788 0 -1 1705
box -2 -3 42 103
use INVX1  INVX1_119
timestamp 1719641852
transform 1 0 764 0 1 1505
box -2 -3 18 103
use INVX1  INVX1_80
timestamp 1719641852
transform 1 0 748 0 1 1505
box -2 -3 18 103
use OAI21X1  OAI21X1_39
timestamp 1719641852
transform 1 0 788 0 -1 1705
box -2 -3 34 103
use BUFX4  BUFX4_23
timestamp 1719641852
transform 1 0 812 0 1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_68
timestamp 1719641852
transform 1 0 780 0 1 1505
box -2 -3 34 103
use FILL  FILL_16_1_1
timestamp 1719641852
transform -1 0 868 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_1_0
timestamp 1719641852
transform -1 0 860 0 -1 1705
box -2 -3 10 103
use OAI21X1  OAI21X1_69
timestamp 1719641852
transform -1 0 852 0 -1 1705
box -2 -3 34 103
use BUFX4  BUFX4_11
timestamp 1719641852
transform 1 0 860 0 1 1505
box -2 -3 34 103
use FILL  FILL_15_1_1
timestamp 1719641852
transform 1 0 852 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_1_0
timestamp 1719641852
transform 1 0 844 0 1 1505
box -2 -3 10 103
use OAI22X1  OAI22X1_30
timestamp 1719641852
transform 1 0 900 0 -1 1705
box -2 -3 42 103
use BUFX4  BUFX4_202
timestamp 1719641852
transform -1 0 900 0 -1 1705
box -2 -3 34 103
use BUFX4  BUFX4_10
timestamp 1719641852
transform 1 0 892 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_16
timestamp 1719641852
transform 1 0 940 0 -1 1705
box -2 -3 26 103
use BUFX4  BUFX4_9
timestamp 1719641852
transform 1 0 924 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_13
timestamp 1719641852
transform -1 0 1012 0 -1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_17
timestamp 1719641852
transform 1 0 964 0 -1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_57
timestamp 1719641852
transform -1 0 1020 0 1 1505
box -2 -3 26 103
use OAI22X1  OAI22X1_31
timestamp 1719641852
transform 1 0 956 0 1 1505
box -2 -3 42 103
use BUFX4  BUFX4_227
timestamp 1719641852
transform 1 0 1036 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_51
timestamp 1719641852
transform -1 0 1036 0 -1 1705
box -2 -3 26 103
use BUFX4  BUFX4_199
timestamp 1719641852
transform -1 0 1052 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_15
timestamp 1719641852
transform 1 0 1068 0 -1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_52
timestamp 1719641852
transform -1 0 1108 0 1 1505
box -2 -3 26 103
use BUFX4  BUFX4_226
timestamp 1719641852
transform 1 0 1052 0 1 1505
box -2 -3 34 103
use INVX2  INVX2_87
timestamp 1719641852
transform 1 0 1180 0 -1 1705
box -2 -3 18 103
use NAND2X1  NAND2X1_233
timestamp 1719641852
transform -1 0 1180 0 -1 1705
box -2 -3 26 103
use INVX8  INVX8_6
timestamp 1719641852
transform 1 0 1116 0 -1 1705
box -2 -3 42 103
use NAND2X1  NAND2X1_54
timestamp 1719641852
transform -1 0 1116 0 -1 1705
box -2 -3 26 103
use INVX1  INVX1_56
timestamp 1719641852
transform -1 0 1188 0 1 1505
box -2 -3 18 103
use INVX1  INVX1_48
timestamp 1719641852
transform -1 0 1172 0 1 1505
box -2 -3 18 103
use NAND2X1  NAND2X1_232
timestamp 1719641852
transform -1 0 1156 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_238
timestamp 1719641852
transform -1 0 1132 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_699
timestamp 1719641852
transform 1 0 1260 0 -1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_9
timestamp 1719641852
transform 1 0 1228 0 -1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_84
timestamp 1719641852
transform 1 0 1196 0 -1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_82
timestamp 1719641852
transform 1 0 1188 0 1 1505
box -2 -3 34 103
use DFFSR  DFFSR_135
timestamp 1719641852
transform -1 0 1396 0 1 1505
box -2 -3 178 103
use NAND2X1  NAND2X1_308
timestamp 1719641852
transform -1 0 1316 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_702
timestamp 1719641852
transform -1 0 1348 0 -1 1705
box -2 -3 34 103
use FILL  FILL_16_2_0
timestamp 1719641852
transform -1 0 1388 0 -1 1705
box -2 -3 10 103
use AOI21X1  AOI21X1_10
timestamp 1719641852
transform 1 0 1348 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_683
timestamp 1719641852
transform -1 0 1428 0 -1 1705
box -2 -3 34 103
use FILL  FILL_16_2_1
timestamp 1719641852
transform -1 0 1396 0 -1 1705
box -2 -3 10 103
use NAND3X1  NAND3X1_78
timestamp 1719641852
transform 1 0 1412 0 1 1505
box -2 -3 34 103
use FILL  FILL_15_2_1
timestamp 1719641852
transform 1 0 1404 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_2_0
timestamp 1719641852
transform 1 0 1396 0 1 1505
box -2 -3 10 103
use OAI21X1  OAI21X1_682
timestamp 1719641852
transform -1 0 1460 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_700
timestamp 1719641852
transform 1 0 1444 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_321
timestamp 1719641852
transform -1 0 1556 0 -1 1705
box -2 -3 26 103
use INVX1  INVX1_151
timestamp 1719641852
transform 1 0 1516 0 -1 1705
box -2 -3 18 103
use OAI21X1  OAI21X1_681
timestamp 1719641852
transform -1 0 1516 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_298
timestamp 1719641852
transform 1 0 1460 0 -1 1705
box -2 -3 26 103
use OR2X2  OR2X2_18
timestamp 1719641852
transform -1 0 1572 0 1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_80
timestamp 1719641852
transform 1 0 1508 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_701
timestamp 1719641852
transform -1 0 1508 0 1 1505
box -2 -3 34 103
use BUFX4  BUFX4_125
timestamp 1719641852
transform -1 0 1620 0 1 1505
box -2 -3 34 103
use INVX1  INVX1_55
timestamp 1719641852
transform -1 0 1588 0 1 1505
box -2 -3 18 103
use DFFSR  DFFSR_168
timestamp 1719641852
transform 1 0 1556 0 -1 1705
box -2 -3 178 103
use DFFSR  DFFSR_156
timestamp 1719641852
transform -1 0 1796 0 1 1505
box -2 -3 178 103
use NOR2X1  NOR2X1_288
timestamp 1719641852
transform 1 0 1796 0 1 1505
box -2 -3 26 103
use AOI22X1  AOI22X1_9
timestamp 1719641852
transform 1 0 1732 0 -1 1705
box -2 -3 42 103
use AOI21X1  AOI21X1_206
timestamp 1719641852
transform 1 0 1772 0 -1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_277
timestamp 1719641852
transform -1 0 1828 0 -1 1705
box -2 -3 26 103
use AOI21X1  AOI21X1_229
timestamp 1719641852
transform -1 0 1852 0 1 1505
box -2 -3 34 103
use INVX2  INVX2_88
timestamp 1719641852
transform 1 0 1828 0 -1 1705
box -2 -3 18 103
use OAI21X1  OAI21X1_593
timestamp 1719641852
transform 1 0 1844 0 -1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_228
timestamp 1719641852
transform -1 0 1884 0 1 1505
box -2 -3 34 103
use FILL  FILL_15_3_0
timestamp 1719641852
transform 1 0 1884 0 1 1505
box -2 -3 10 103
use FILL  FILL_16_3_0
timestamp 1719641852
transform 1 0 1876 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_3_1
timestamp 1719641852
transform 1 0 1884 0 -1 1705
box -2 -3 10 103
use FILL  FILL_15_3_1
timestamp 1719641852
transform 1 0 1892 0 1 1505
box -2 -3 10 103
use BUFX4  BUFX4_203
timestamp 1719641852
transform 1 0 1900 0 1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_204
timestamp 1719641852
transform 1 0 1892 0 -1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_209
timestamp 1719641852
transform -1 0 1996 0 -1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_279
timestamp 1719641852
transform 1 0 1940 0 -1 1705
box -2 -3 26 103
use INVX2  INVX2_121
timestamp 1719641852
transform 1 0 1924 0 -1 1705
box -2 -3 18 103
use DFFSR  DFFSR_167
timestamp 1719641852
transform -1 0 2108 0 1 1505
box -2 -3 178 103
use DFFSR  DFFSR_171
timestamp 1719641852
transform -1 0 2284 0 1 1505
box -2 -3 178 103
use OAI21X1  OAI21X1_595
timestamp 1719641852
transform 1 0 1996 0 -1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_207
timestamp 1719641852
transform -1 0 2060 0 -1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_334
timestamp 1719641852
transform -1 0 2084 0 -1 1705
box -2 -3 26 103
use AOI22X1  AOI22X1_16
timestamp 1719641852
transform 1 0 2084 0 -1 1705
box -2 -3 42 103
use INVX2  INVX2_129
timestamp 1719641852
transform 1 0 2124 0 -1 1705
box -2 -3 18 103
use DFFSR  DFFSR_231
timestamp 1719641852
transform -1 0 2316 0 -1 1705
box -2 -3 178 103
use INVX1  INVX1_46
timestamp 1719641852
transform -1 0 2300 0 1 1505
box -2 -3 18 103
use BUFX4  BUFX4_39
timestamp 1719641852
transform 1 0 2300 0 1 1505
box -2 -3 34 103
use FILL  FILL_15_4_0
timestamp 1719641852
transform -1 0 2340 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_4_1
timestamp 1719641852
transform -1 0 2348 0 1 1505
box -2 -3 10 103
use DFFSR  DFFSR_200
timestamp 1719641852
transform -1 0 2524 0 1 1505
box -2 -3 178 103
use OR2X2  OR2X2_15
timestamp 1719641852
transform 1 0 2316 0 -1 1705
box -2 -3 34 103
use FILL  FILL_16_4_0
timestamp 1719641852
transform -1 0 2356 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_4_1
timestamp 1719641852
transform -1 0 2364 0 -1 1705
box -2 -3 10 103
use NOR2X1  NOR2X1_247
timestamp 1719641852
transform -1 0 2548 0 1 1505
box -2 -3 26 103
use DFFSR  DFFSR_215
timestamp 1719641852
transform -1 0 2540 0 -1 1705
box -2 -3 178 103
use OAI21X1  OAI21X1_472
timestamp 1719641852
transform -1 0 2636 0 -1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_165
timestamp 1719641852
transform 1 0 2572 0 -1 1705
box -2 -3 34 103
use INVX2  INVX2_114
timestamp 1719641852
transform -1 0 2572 0 -1 1705
box -2 -3 18 103
use INVX2  INVX2_91
timestamp 1719641852
transform 1 0 2540 0 -1 1705
box -2 -3 18 103
use BUFX4  BUFX4_49
timestamp 1719641852
transform -1 0 2644 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_474
timestamp 1719641852
transform -1 0 2612 0 1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_166
timestamp 1719641852
transform -1 0 2580 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_362
timestamp 1719641852
transform 1 0 2716 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_361
timestamp 1719641852
transform -1 0 2716 0 -1 1705
box -2 -3 34 103
use INVX2  INVX2_162
timestamp 1719641852
transform 1 0 2668 0 -1 1705
box -2 -3 18 103
use BUFX4  BUFX4_232
timestamp 1719641852
transform 1 0 2636 0 -1 1705
box -2 -3 34 103
use INVX2  INVX2_128
timestamp 1719641852
transform 1 0 2660 0 1 1505
box -2 -3 18 103
use INVX2  INVX2_158
timestamp 1719641852
transform 1 0 2644 0 1 1505
box -2 -3 18 103
use DFFSR  DFFSR_233
timestamp 1719641852
transform -1 0 2852 0 1 1505
box -2 -3 178 103
use OAI21X1  OAI21X1_365
timestamp 1719641852
transform -1 0 2884 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_364
timestamp 1719641852
transform 1 0 2884 0 1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_112
timestamp 1719641852
transform -1 0 2780 0 -1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_119
timestamp 1719641852
transform -1 0 2812 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_371
timestamp 1719641852
transform -1 0 2844 0 -1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_215
timestamp 1719641852
transform 1 0 2844 0 -1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_212
timestamp 1719641852
transform -1 0 2892 0 -1 1705
box -2 -3 26 103
use FILL  FILL_16_5_0
timestamp 1719641852
transform 1 0 2892 0 -1 1705
box -2 -3 10 103
use AOI21X1  AOI21X1_140
timestamp 1719641852
transform 1 0 2908 0 -1 1705
box -2 -3 34 103
use FILL  FILL_16_5_1
timestamp 1719641852
transform 1 0 2900 0 -1 1705
box -2 -3 10 103
use BUFX4  BUFX4_50
timestamp 1719641852
transform 1 0 2932 0 1 1505
box -2 -3 34 103
use FILL  FILL_15_5_1
timestamp 1719641852
transform 1 0 2924 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_5_0
timestamp 1719641852
transform 1 0 2916 0 1 1505
box -2 -3 10 103
use INVX1  INVX1_128
timestamp 1719641852
transform -1 0 2988 0 -1 1705
box -2 -3 18 103
use OAI21X1  OAI21X1_424
timestamp 1719641852
transform -1 0 2972 0 -1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_251
timestamp 1719641852
transform -1 0 2996 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_228
timestamp 1719641852
transform -1 0 3012 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_747
timestamp 1719641852
transform -1 0 3028 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_213
timestamp 1719641852
transform -1 0 3068 0 -1 1705
box -2 -3 26 103
use BUFX4  BUFX4_230
timestamp 1719641852
transform -1 0 3044 0 -1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_327
timestamp 1719641852
transform -1 0 3052 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_223
timestamp 1719641852
transform 1 0 3068 0 -1 1705
box -2 -3 26 103
use AOI21X1  AOI21X1_136
timestamp 1719641852
transform 1 0 3076 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_226
timestamp 1719641852
transform -1 0 3076 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_227
timestamp 1719641852
transform -1 0 3140 0 -1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_217
timestamp 1719641852
transform -1 0 3116 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_417
timestamp 1719641852
transform -1 0 3140 0 1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_88
timestamp 1719641852
transform -1 0 3172 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_215
timestamp 1719641852
transform -1 0 3188 0 1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_195
timestamp 1719641852
transform -1 0 3164 0 1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_86
timestamp 1719641852
transform -1 0 3244 0 -1 1705
box -2 -3 34 103
use INVX8  INVX8_14
timestamp 1719641852
transform 1 0 3172 0 -1 1705
box -2 -3 42 103
use NAND2X1  NAND2X1_329
timestamp 1719641852
transform -1 0 3236 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_220
timestamp 1719641852
transform -1 0 3212 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_185
timestamp 1719641852
transform -1 0 3268 0 -1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_194
timestamp 1719641852
transform 1 0 3260 0 1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_198
timestamp 1719641852
transform 1 0 3236 0 1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_183
timestamp 1719641852
transform 1 0 3292 0 -1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_191
timestamp 1719641852
transform 1 0 3268 0 -1 1705
box -2 -3 26 103
use AOI22X1  AOI22X1_46
timestamp 1719641852
transform 1 0 3284 0 1 1505
box -2 -3 42 103
use AOI21X1  AOI21X1_79
timestamp 1719641852
transform -1 0 3372 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_181
timestamp 1719641852
transform 1 0 3316 0 -1 1705
box -2 -3 26 103
use AOI21X1  AOI21X1_67
timestamp 1719641852
transform -1 0 3356 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_105
timestamp 1719641852
transform 1 0 3396 0 -1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_143
timestamp 1719641852
transform 1 0 3372 0 -1 1705
box -2 -3 26 103
use AOI22X1  AOI22X1_50
timestamp 1719641852
transform 1 0 3396 0 1 1505
box -2 -3 42 103
use AOI22X1  AOI22X1_41
timestamp 1719641852
transform 1 0 3356 0 1 1505
box -2 -3 42 103
use NOR2X1  NOR2X1_106
timestamp 1719641852
transform 1 0 3436 0 -1 1705
box -2 -3 26 103
use FILL  FILL_16_6_1
timestamp 1719641852
transform 1 0 3428 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_6_0
timestamp 1719641852
transform 1 0 3420 0 -1 1705
box -2 -3 10 103
use FILL  FILL_15_6_0
timestamp 1719641852
transform 1 0 3436 0 1 1505
box -2 -3 10 103
use OAI21X1  OAI21X1_223
timestamp 1719641852
transform 1 0 3460 0 -1 1705
box -2 -3 34 103
use AOI22X1  AOI22X1_54
timestamp 1719641852
transform 1 0 3452 0 1 1505
box -2 -3 42 103
use FILL  FILL_15_6_1
timestamp 1719641852
transform 1 0 3444 0 1 1505
box -2 -3 10 103
use OAI21X1  OAI21X1_248
timestamp 1719641852
transform 1 0 3516 0 -1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_142
timestamp 1719641852
transform 1 0 3492 0 -1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_199
timestamp 1719641852
transform 1 0 3524 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_297
timestamp 1719641852
transform -1 0 3524 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_132
timestamp 1719641852
transform 1 0 3572 0 -1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_131
timestamp 1719641852
transform 1 0 3548 0 -1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_186
timestamp 1719641852
transform 1 0 3564 0 1 1505
box -2 -3 26 103
use INVX1  INVX1_109
timestamp 1719641852
transform 1 0 3548 0 1 1505
box -2 -3 18 103
use OAI21X1  OAI21X1_242
timestamp 1719641852
transform 1 0 3596 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_110
timestamp 1719641852
transform 1 0 3620 0 1 1505
box -2 -3 18 103
use OAI21X1  OAI21X1_303
timestamp 1719641852
transform -1 0 3620 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_107
timestamp 1719641852
transform 1 0 3652 0 -1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_108
timestamp 1719641852
transform 1 0 3628 0 -1 1705
box -2 -3 26 103
use BUFX4  BUFX4_215
timestamp 1719641852
transform -1 0 3692 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_185
timestamp 1719641852
transform -1 0 3660 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_224
timestamp 1719641852
transform 1 0 3676 0 -1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_127
timestamp 1719641852
transform -1 0 3724 0 1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_129
timestamp 1719641852
transform -1 0 3740 0 -1 1705
box -2 -3 34 103
use BUFX4  BUFX4_237
timestamp 1719641852
transform -1 0 3756 0 1 1505
box -2 -3 34 103
use NAND3X1  NAND3X1_131
timestamp 1719641852
transform -1 0 3772 0 -1 1705
box -2 -3 34 103
use FILL  FILL_16_2
timestamp 1719641852
transform 1 0 3764 0 1 1505
box -2 -3 10 103
use FILL  FILL_16_1
timestamp 1719641852
transform 1 0 3756 0 1 1505
box -2 -3 10 103
use FILL  FILL_17_1
timestamp 1719641852
transform -1 0 3780 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_3
timestamp 1719641852
transform 1 0 3772 0 1 1505
box -2 -3 10 103
use BUFX2  BUFX2_47
timestamp 1719641852
transform -1 0 28 0 1 1705
box -2 -3 26 103
use DFFSR  DFFSR_76
timestamp 1719641852
transform -1 0 204 0 1 1705
box -2 -3 178 103
use CLKBUF1  CLKBUF1_47
timestamp 1719641852
transform -1 0 276 0 1 1705
box -2 -3 74 103
use NOR2X1  NOR2X1_35
timestamp 1719641852
transform 1 0 276 0 1 1705
box -2 -3 26 103
use NAND3X1  NAND3X1_105
timestamp 1719641852
transform 1 0 300 0 1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_36
timestamp 1719641852
transform -1 0 356 0 1 1705
box -2 -3 26 103
use FILL  FILL_17_0_0
timestamp 1719641852
transform -1 0 364 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_0_1
timestamp 1719641852
transform -1 0 372 0 1 1705
box -2 -3 10 103
use NOR2X1  NOR2X1_38
timestamp 1719641852
transform -1 0 396 0 1 1705
box -2 -3 26 103
use OR2X2  OR2X2_2
timestamp 1719641852
transform -1 0 428 0 1 1705
box -2 -3 34 103
use INVX2  INVX2_28
timestamp 1719641852
transform 1 0 428 0 1 1705
box -2 -3 18 103
use OAI21X1  OAI21X1_95
timestamp 1719641852
transform 1 0 444 0 1 1705
box -2 -3 34 103
use INVX2  INVX2_23
timestamp 1719641852
transform -1 0 492 0 1 1705
box -2 -3 18 103
use OAI21X1  OAI21X1_105
timestamp 1719641852
transform 1 0 492 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_104
timestamp 1719641852
transform 1 0 524 0 1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_56
timestamp 1719641852
transform 1 0 556 0 1 1705
box -2 -3 34 103
use BUFX4  BUFX4_94
timestamp 1719641852
transform 1 0 588 0 1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_51
timestamp 1719641852
transform 1 0 620 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_94
timestamp 1719641852
transform -1 0 684 0 1 1705
box -2 -3 34 103
use AND2X2  AND2X2_3
timestamp 1719641852
transform 1 0 684 0 1 1705
box -2 -3 34 103
use INVX8  INVX8_4
timestamp 1719641852
transform -1 0 756 0 1 1705
box -2 -3 42 103
use OAI22X1  OAI22X1_32
timestamp 1719641852
transform -1 0 796 0 1 1705
box -2 -3 42 103
use NAND3X1  NAND3X1_22
timestamp 1719641852
transform 1 0 796 0 1 1705
box -2 -3 34 103
use OAI22X1  OAI22X1_22
timestamp 1719641852
transform 1 0 828 0 1 1705
box -2 -3 42 103
use FILL  FILL_17_1_0
timestamp 1719641852
transform -1 0 876 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_1_1
timestamp 1719641852
transform -1 0 884 0 1 1705
box -2 -3 10 103
use NOR2X1  NOR2X1_12
timestamp 1719641852
transform -1 0 908 0 1 1705
box -2 -3 26 103
use OAI22X1  OAI22X1_21
timestamp 1719641852
transform 1 0 908 0 1 1705
box -2 -3 42 103
use BUFX4  BUFX4_76
timestamp 1719641852
transform -1 0 980 0 1 1705
box -2 -3 34 103
use INVX1  INVX1_47
timestamp 1719641852
transform -1 0 996 0 1 1705
box -2 -3 18 103
use OAI22X1  OAI22X1_23
timestamp 1719641852
transform 1 0 996 0 1 1705
box -2 -3 42 103
use BUFX4  BUFX4_77
timestamp 1719641852
transform 1 0 1036 0 1 1705
box -2 -3 34 103
use DFFSR  DFFSR_128
timestamp 1719641852
transform -1 0 1244 0 1 1705
box -2 -3 178 103
use NAND2X1  NAND2X1_48
timestamp 1719641852
transform -1 0 1268 0 1 1705
box -2 -3 26 103
use DFFSR  DFFSR_218
timestamp 1719641852
transform -1 0 1444 0 1 1705
box -2 -3 178 103
use FILL  FILL_17_2_0
timestamp 1719641852
transform 1 0 1444 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_2_1
timestamp 1719641852
transform 1 0 1452 0 1 1705
box -2 -3 10 103
use NAND2X1  NAND2X1_297
timestamp 1719641852
transform 1 0 1460 0 1 1705
box -2 -3 26 103
use INVX2  INVX2_119
timestamp 1719641852
transform 1 0 1484 0 1 1705
box -2 -3 18 103
use NAND2X1  NAND2X1_50
timestamp 1719641852
transform -1 0 1524 0 1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_321
timestamp 1719641852
transform -1 0 1548 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_679
timestamp 1719641852
transform -1 0 1580 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_723
timestamp 1719641852
transform -1 0 1612 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_680
timestamp 1719641852
transform 1 0 1612 0 1 1705
box -2 -3 34 103
use CLKBUF1  CLKBUF1_50
timestamp 1719641852
transform 1 0 1644 0 1 1705
box -2 -3 74 103
use BUFX4  BUFX4_31
timestamp 1719641852
transform -1 0 1748 0 1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_205
timestamp 1719641852
transform 1 0 1748 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_594
timestamp 1719641852
transform -1 0 1812 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_596
timestamp 1719641852
transform -1 0 1844 0 1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_208
timestamp 1719641852
transform 1 0 1844 0 1 1705
box -2 -3 34 103
use FILL  FILL_17_3_0
timestamp 1719641852
transform -1 0 1884 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_3_1
timestamp 1719641852
transform -1 0 1892 0 1 1705
box -2 -3 10 103
use NAND2X1  NAND2X1_265
timestamp 1719641852
transform -1 0 1916 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_772
timestamp 1719641852
transform 1 0 1916 0 1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_261
timestamp 1719641852
transform -1 0 1980 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_266
timestamp 1719641852
transform 1 0 1980 0 1 1705
box -2 -3 26 103
use AOI21X1  AOI21X1_262
timestamp 1719641852
transform 1 0 2004 0 1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_263
timestamp 1719641852
transform 1 0 2036 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_773
timestamp 1719641852
transform -1 0 2100 0 1 1705
box -2 -3 34 103
use INVX2  INVX2_118
timestamp 1719641852
transform -1 0 2116 0 1 1705
box -2 -3 18 103
use NOR2X1  NOR2X1_278
timestamp 1719641852
transform -1 0 2140 0 1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_276
timestamp 1719641852
transform 1 0 2140 0 1 1705
box -2 -3 26 103
use INVX8  INVX8_19
timestamp 1719641852
transform -1 0 2204 0 1 1705
box -2 -3 42 103
use NOR2X1  NOR2X1_214
timestamp 1719641852
transform 1 0 2204 0 1 1705
box -2 -3 26 103
use AOI21X1  AOI21X1_118
timestamp 1719641852
transform -1 0 2260 0 1 1705
box -2 -3 34 103
use DFFSR  DFFSR_230
timestamp 1719641852
transform -1 0 2436 0 1 1705
box -2 -3 178 103
use FILL  FILL_17_4_0
timestamp 1719641852
transform -1 0 2444 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_4_1
timestamp 1719641852
transform -1 0 2452 0 1 1705
box -2 -3 10 103
use OAI21X1  OAI21X1_411
timestamp 1719641852
transform -1 0 2484 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_415
timestamp 1719641852
transform -1 0 2516 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_363
timestamp 1719641852
transform -1 0 2548 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_427
timestamp 1719641852
transform -1 0 2580 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_423
timestamp 1719641852
transform -1 0 2612 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_473
timestamp 1719641852
transform -1 0 2644 0 1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_135
timestamp 1719641852
transform -1 0 2676 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_412
timestamp 1719641852
transform -1 0 2708 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_748
timestamp 1719641852
transform -1 0 2740 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_373
timestamp 1719641852
transform 1 0 2740 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_374
timestamp 1719641852
transform 1 0 2772 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_370
timestamp 1719641852
transform -1 0 2836 0 1 1705
box -2 -3 34 103
use BUFX4  BUFX4_244
timestamp 1719641852
transform -1 0 2868 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_368
timestamp 1719641852
transform 1 0 2868 0 1 1705
box -2 -3 34 103
use FILL  FILL_17_5_0
timestamp 1719641852
transform -1 0 2908 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_5_1
timestamp 1719641852
transform -1 0 2916 0 1 1705
box -2 -3 10 103
use AOI21X1  AOI21X1_116
timestamp 1719641852
transform -1 0 2948 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_221
timestamp 1719641852
transform -1 0 2972 0 1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_225
timestamp 1719641852
transform 1 0 2972 0 1 1705
box -2 -3 26 103
use BUFX4  BUFX4_52
timestamp 1719641852
transform -1 0 3028 0 1 1705
box -2 -3 34 103
use INVX8  INVX8_15
timestamp 1719641852
transform 1 0 3028 0 1 1705
box -2 -3 42 103
use INVX1  INVX1_127
timestamp 1719641852
transform -1 0 3084 0 1 1705
box -2 -3 18 103
use AOI22X1  AOI22X1_57
timestamp 1719641852
transform -1 0 3124 0 1 1705
box -2 -3 42 103
use OAI21X1  OAI21X1_304
timestamp 1719641852
transform 1 0 3124 0 1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_204
timestamp 1719641852
transform 1 0 3156 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_187
timestamp 1719641852
transform -1 0 3212 0 1 1705
box -2 -3 26 103
use AOI22X1  AOI22X1_55
timestamp 1719641852
transform 1 0 3212 0 1 1705
box -2 -3 42 103
use NAND2X1  NAND2X1_186
timestamp 1719641852
transform -1 0 3276 0 1 1705
box -2 -3 26 103
use INVX1  INVX1_114
timestamp 1719641852
transform -1 0 3292 0 1 1705
box -2 -3 18 103
use AOI21X1  AOI21X1_80
timestamp 1719641852
transform 1 0 3292 0 1 1705
box -2 -3 34 103
use AOI22X1  AOI22X1_52
timestamp 1719641852
transform -1 0 3364 0 1 1705
box -2 -3 42 103
use NAND2X1  NAND2X1_180
timestamp 1719641852
transform -1 0 3388 0 1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_182
timestamp 1719641852
transform 1 0 3388 0 1 1705
box -2 -3 26 103
use FILL  FILL_17_6_0
timestamp 1719641852
transform -1 0 3420 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_6_1
timestamp 1719641852
transform -1 0 3428 0 1 1705
box -2 -3 10 103
use BUFX4  BUFX4_174
timestamp 1719641852
transform -1 0 3460 0 1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_134
timestamp 1719641852
transform 1 0 3460 0 1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_133
timestamp 1719641852
transform 1 0 3484 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_243
timestamp 1719641852
transform 1 0 3508 0 1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_151
timestamp 1719641852
transform -1 0 3572 0 1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_153
timestamp 1719641852
transform -1 0 3604 0 1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_145
timestamp 1719641852
transform -1 0 3636 0 1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_146
timestamp 1719641852
transform 1 0 3636 0 1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_147
timestamp 1719641852
transform -1 0 3700 0 1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_154
timestamp 1719641852
transform -1 0 3732 0 1 1705
box -2 -3 34 103
use INVX2  INVX2_47
timestamp 1719641852
transform 1 0 3732 0 1 1705
box -2 -3 18 103
use NAND3X1  NAND3X1_132
timestamp 1719641852
transform -1 0 3780 0 1 1705
box -2 -3 34 103
use INVX8  INVX8_3
timestamp 1719641852
transform -1 0 44 0 -1 1905
box -2 -3 42 103
use DFFSR  DFFSR_46
timestamp 1719641852
transform -1 0 220 0 -1 1905
box -2 -3 178 103
use INVX2  INVX2_4
timestamp 1719641852
transform 1 0 220 0 -1 1905
box -2 -3 18 103
use DFFSR  DFFSR_55
timestamp 1719641852
transform 1 0 236 0 -1 1905
box -2 -3 178 103
use FILL  FILL_18_0_0
timestamp 1719641852
transform -1 0 420 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_0_1
timestamp 1719641852
transform -1 0 428 0 -1 1905
box -2 -3 10 103
use BUFX4  BUFX4_141
timestamp 1719641852
transform -1 0 460 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_36
timestamp 1719641852
transform 1 0 460 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_43
timestamp 1719641852
transform 1 0 492 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_73
timestamp 1719641852
transform -1 0 556 0 -1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_20
timestamp 1719641852
transform 1 0 556 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_35
timestamp 1719641852
transform 1 0 588 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_45
timestamp 1719641852
transform 1 0 620 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_17
timestamp 1719641852
transform 1 0 652 0 -1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_40
timestamp 1719641852
transform 1 0 676 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_65
timestamp 1719641852
transform 1 0 708 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_170
timestamp 1719641852
transform 1 0 740 0 -1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_298
timestamp 1719641852
transform -1 0 796 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_103
timestamp 1719641852
transform -1 0 820 0 -1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_56
timestamp 1719641852
transform -1 0 844 0 -1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_49
timestamp 1719641852
transform -1 0 868 0 -1 1905
box -2 -3 26 103
use FILL  FILL_18_1_0
timestamp 1719641852
transform -1 0 876 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_1_1
timestamp 1719641852
transform -1 0 884 0 -1 1905
box -2 -3 10 103
use NAND3X1  NAND3X1_83
timestamp 1719641852
transform -1 0 916 0 -1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_13
timestamp 1719641852
transform -1 0 948 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_55
timestamp 1719641852
transform -1 0 972 0 -1 1905
box -2 -3 26 103
use NAND3X1  NAND3X1_79
timestamp 1719641852
transform -1 0 1004 0 -1 1905
box -2 -3 34 103
use NOR3X1  NOR3X1_1
timestamp 1719641852
transform -1 0 1068 0 -1 1905
box -2 -3 66 103
use BUFX4  BUFX4_189
timestamp 1719641852
transform -1 0 1100 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_34
timestamp 1719641852
transform 1 0 1100 0 -1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_126
timestamp 1719641852
transform 1 0 1124 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_35
timestamp 1719641852
transform 1 0 1156 0 -1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_19
timestamp 1719641852
transform -1 0 1204 0 -1 1905
box -2 -3 26 103
use INVX1  INVX1_132
timestamp 1719641852
transform 1 0 1204 0 -1 1905
box -2 -3 18 103
use NAND2X1  NAND2X1_63
timestamp 1719641852
transform -1 0 1244 0 -1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_725
timestamp 1719641852
transform -1 0 1276 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_724
timestamp 1719641852
transform -1 0 1308 0 -1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_234
timestamp 1719641852
transform -1 0 1332 0 -1 1905
box -2 -3 26 103
use CLKBUF1  CLKBUF1_19
timestamp 1719641852
transform 1 0 1332 0 -1 1905
box -2 -3 74 103
use FILL  FILL_18_2_0
timestamp 1719641852
transform 1 0 1404 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_2_1
timestamp 1719641852
transform 1 0 1412 0 -1 1905
box -2 -3 10 103
use NAND3X1  NAND3X1_81
timestamp 1719641852
transform 1 0 1420 0 -1 1905
box -2 -3 34 103
use INVX8  INVX8_18
timestamp 1719641852
transform -1 0 1492 0 -1 1905
box -2 -3 42 103
use INVX4  INVX4_6
timestamp 1719641852
transform -1 0 1516 0 -1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_296
timestamp 1719641852
transform 1 0 1516 0 -1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_319
timestamp 1719641852
transform 1 0 1540 0 -1 1905
box -2 -3 26 103
use INVX1  INVX1_150
timestamp 1719641852
transform -1 0 1580 0 -1 1905
box -2 -3 18 103
use NAND2X1  NAND2X1_278
timestamp 1719641852
transform 1 0 1580 0 -1 1905
box -2 -3 26 103
use AOI22X1  AOI22X1_7
timestamp 1719641852
transform -1 0 1644 0 -1 1905
box -2 -3 42 103
use OAI21X1  OAI21X1_675
timestamp 1719641852
transform -1 0 1676 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_279
timestamp 1719641852
transform 1 0 1676 0 -1 1905
box -2 -3 26 103
use DFFSR  DFFSR_199
timestamp 1719641852
transform -1 0 1876 0 -1 1905
box -2 -3 178 103
use FILL  FILL_18_3_0
timestamp 1719641852
transform 1 0 1876 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_3_1
timestamp 1719641852
transform 1 0 1884 0 -1 1905
box -2 -3 10 103
use OAI21X1  OAI21X1_475
timestamp 1719641852
transform 1 0 1892 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_480
timestamp 1719641852
transform -1 0 1956 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_479
timestamp 1719641852
transform -1 0 1988 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_478
timestamp 1719641852
transform -1 0 2020 0 -1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_167
timestamp 1719641852
transform 1 0 2020 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_477
timestamp 1719641852
transform -1 0 2084 0 -1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_248
timestamp 1719641852
transform 1 0 2084 0 -1 1905
box -2 -3 26 103
use DFFSR  DFFSR_201
timestamp 1719641852
transform 1 0 2108 0 -1 1905
box -2 -3 178 103
use INVX2  INVX2_120
timestamp 1719641852
transform 1 0 2284 0 -1 1905
box -2 -3 18 103
use OAI21X1  OAI21X1_471
timestamp 1719641852
transform 1 0 2300 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_241
timestamp 1719641852
transform 1 0 2332 0 -1 1905
box -2 -3 26 103
use AOI22X1  AOI22X1_11
timestamp 1719641852
transform -1 0 2396 0 -1 1905
box -2 -3 42 103
use FILL  FILL_18_4_0
timestamp 1719641852
transform -1 0 2404 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_4_1
timestamp 1719641852
transform -1 0 2412 0 -1 1905
box -2 -3 10 103
use NOR2X1  NOR2X1_246
timestamp 1719641852
transform -1 0 2436 0 -1 1905
box -2 -3 26 103
use AOI21X1  AOI21X1_164
timestamp 1719641852
transform -1 0 2468 0 -1 1905
box -2 -3 34 103
use INVX2  INVX2_160
timestamp 1719641852
transform 1 0 2468 0 -1 1905
box -2 -3 18 103
use OAI21X1  OAI21X1_414
timestamp 1719641852
transform -1 0 2516 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_476
timestamp 1719641852
transform 1 0 2516 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_426
timestamp 1719641852
transform 1 0 2548 0 -1 1905
box -2 -3 34 103
use DFFSR  DFFSR_203
timestamp 1719641852
transform 1 0 2580 0 -1 1905
box -2 -3 178 103
use NAND2X1  NAND2X1_252
timestamp 1719641852
transform 1 0 2756 0 -1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_468
timestamp 1719641852
transform 1 0 2780 0 -1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_163
timestamp 1719641852
transform 1 0 2812 0 -1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_245
timestamp 1719641852
transform 1 0 2844 0 -1 1905
box -2 -3 26 103
use BUFX4  BUFX4_150
timestamp 1719641852
transform -1 0 2900 0 -1 1905
box -2 -3 34 103
use FILL  FILL_18_5_0
timestamp 1719641852
transform 1 0 2900 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_5_1
timestamp 1719641852
transform 1 0 2908 0 -1 1905
box -2 -3 10 103
use INVX1  INVX1_129
timestamp 1719641852
transform 1 0 2916 0 -1 1905
box -2 -3 18 103
use NAND2X1  NAND2X1_246
timestamp 1719641852
transform 1 0 2932 0 -1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_228
timestamp 1719641852
transform -1 0 2980 0 -1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_218
timestamp 1719641852
transform -1 0 3004 0 -1 1905
box -2 -3 26 103
use BUFX4  BUFX4_241
timestamp 1719641852
transform -1 0 3036 0 -1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_330
timestamp 1719641852
transform 1 0 3036 0 -1 1905
box -2 -3 26 103
use OR2X2  OR2X2_21
timestamp 1719641852
transform -1 0 3092 0 -1 1905
box -2 -3 34 103
use BUFX4  BUFX4_59
timestamp 1719641852
transform -1 0 3124 0 -1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_205
timestamp 1719641852
transform -1 0 3156 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_306
timestamp 1719641852
transform 1 0 3156 0 -1 1905
box -2 -3 34 103
use AOI22X1  AOI22X1_56
timestamp 1719641852
transform -1 0 3228 0 -1 1905
box -2 -3 42 103
use NOR2X1  NOR2X1_192
timestamp 1719641852
transform -1 0 3252 0 -1 1905
box -2 -3 26 103
use AOI21X1  AOI21X1_92
timestamp 1719641852
transform -1 0 3284 0 -1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_90
timestamp 1719641852
transform -1 0 3316 0 -1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_87
timestamp 1719641852
transform -1 0 3348 0 -1 1905
box -2 -3 34 103
use BUFX4  BUFX4_156
timestamp 1719641852
transform -1 0 3380 0 -1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_130
timestamp 1719641852
transform 1 0 3380 0 -1 1905
box -2 -3 26 103
use FILL  FILL_18_6_0
timestamp 1719641852
transform 1 0 3404 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_6_1
timestamp 1719641852
transform 1 0 3412 0 -1 1905
box -2 -3 10 103
use OAI21X1  OAI21X1_241
timestamp 1719641852
transform 1 0 3420 0 -1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_144
timestamp 1719641852
transform 1 0 3452 0 -1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_145
timestamp 1719641852
transform 1 0 3476 0 -1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_249
timestamp 1719641852
transform 1 0 3500 0 -1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_127
timestamp 1719641852
transform 1 0 3532 0 -1 1905
box -2 -3 26 103
use NAND3X1  NAND3X1_152
timestamp 1719641852
transform -1 0 3588 0 -1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_128
timestamp 1719641852
transform 1 0 3588 0 -1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_240
timestamp 1719641852
transform 1 0 3612 0 -1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_144
timestamp 1719641852
transform -1 0 3676 0 -1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_130
timestamp 1719641852
transform -1 0 3708 0 -1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_123
timestamp 1719641852
transform -1 0 3740 0 -1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_116
timestamp 1719641852
transform -1 0 3772 0 -1 1905
box -2 -3 34 103
use FILL  FILL_19_1
timestamp 1719641852
transform -1 0 3780 0 -1 1905
box -2 -3 10 103
use BUFX2  BUFX2_14
timestamp 1719641852
transform -1 0 28 0 1 1905
box -2 -3 26 103
use BUFX2  BUFX2_44
timestamp 1719641852
transform -1 0 52 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_138
timestamp 1719641852
transform 1 0 52 0 1 1905
box -2 -3 34 103
use DFFSR  DFFSR_12
timestamp 1719641852
transform -1 0 260 0 1 1905
box -2 -3 178 103
use OAI21X1  OAI21X1_136
timestamp 1719641852
transform 1 0 260 0 1 1905
box -2 -3 34 103
use INVX2  INVX2_6
timestamp 1719641852
transform 1 0 292 0 1 1905
box -2 -3 18 103
use BUFX4  BUFX4_91
timestamp 1719641852
transform -1 0 340 0 1 1905
box -2 -3 34 103
use FILL  FILL_19_0_0
timestamp 1719641852
transform 1 0 340 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_0_1
timestamp 1719641852
transform 1 0 348 0 1 1905
box -2 -3 10 103
use INVX2  INVX2_2
timestamp 1719641852
transform 1 0 356 0 1 1905
box -2 -3 18 103
use DFFSR  DFFSR_10
timestamp 1719641852
transform -1 0 548 0 1 1905
box -2 -3 178 103
use OAI21X1  OAI21X1_74
timestamp 1719641852
transform -1 0 580 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_44
timestamp 1719641852
transform 1 0 580 0 1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_24
timestamp 1719641852
transform 1 0 612 0 1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_23
timestamp 1719641852
transform 1 0 644 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_41
timestamp 1719641852
transform -1 0 708 0 1 1905
box -2 -3 34 103
use INVX1  INVX1_17
timestamp 1719641852
transform -1 0 724 0 1 1905
box -2 -3 18 103
use DFFSR  DFFSR_73
timestamp 1719641852
transform -1 0 900 0 1 1905
box -2 -3 178 103
use FILL  FILL_19_1_0
timestamp 1719641852
transform -1 0 908 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_1_1
timestamp 1719641852
transform -1 0 916 0 1 1905
box -2 -3 10 103
use OAI21X1  OAI21X1_67
timestamp 1719641852
transform -1 0 948 0 1 1905
box -2 -3 34 103
use INVX1  INVX1_18
timestamp 1719641852
transform -1 0 964 0 1 1905
box -2 -3 18 103
use BUFX4  BUFX4_20
timestamp 1719641852
transform -1 0 996 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_181
timestamp 1719641852
transform -1 0 1028 0 1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_2
timestamp 1719641852
transform -1 0 1060 0 1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_50
timestamp 1719641852
transform 1 0 1060 0 1 1905
box -2 -3 34 103
use INVX4  INVX4_1
timestamp 1719641852
transform 1 0 1092 0 1 1905
box -2 -3 26 103
use NAND3X1  NAND3X1_35
timestamp 1719641852
transform 1 0 1116 0 1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_75
timestamp 1719641852
transform -1 0 1180 0 1 1905
box -2 -3 34 103
use INVX2  INVX2_39
timestamp 1719641852
transform -1 0 1196 0 1 1905
box -2 -3 18 103
use DFFSR  DFFSR_119
timestamp 1719641852
transform 1 0 1196 0 1 1905
box -2 -3 178 103
use FILL  FILL_19_2_0
timestamp 1719641852
transform 1 0 1372 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_2_1
timestamp 1719641852
transform 1 0 1380 0 1 1905
box -2 -3 10 103
use INVX2  INVX2_117
timestamp 1719641852
transform 1 0 1388 0 1 1905
box -2 -3 18 103
use NAND2X1  NAND2X1_320
timestamp 1719641852
transform 1 0 1404 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_722
timestamp 1719641852
transform -1 0 1460 0 1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_89
timestamp 1719641852
transform 1 0 1460 0 1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_22
timestamp 1719641852
transform -1 0 1516 0 1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_20
timestamp 1719641852
transform -1 0 1540 0 1 1905
box -2 -3 26 103
use INVX1  INVX1_40
timestamp 1719641852
transform -1 0 1556 0 1 1905
box -2 -3 18 103
use OAI21X1  OAI21X1_636
timestamp 1719641852
transform 1 0 1556 0 1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_234
timestamp 1719641852
transform 1 0 1588 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_720
timestamp 1719641852
transform 1 0 1620 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_719
timestamp 1719641852
transform -1 0 1684 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_266
timestamp 1719641852
transform 1 0 1684 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_677
timestamp 1719641852
transform 1 0 1716 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_676
timestamp 1719641852
transform 1 0 1748 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_638
timestamp 1719641852
transform 1 0 1780 0 1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_237
timestamp 1719641852
transform 1 0 1812 0 1 1905
box -2 -3 34 103
use BUFX4  BUFX4_209
timestamp 1719641852
transform 1 0 1844 0 1 1905
box -2 -3 34 103
use FILL  FILL_19_3_0
timestamp 1719641852
transform 1 0 1876 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_3_1
timestamp 1719641852
transform 1 0 1884 0 1 1905
box -2 -3 10 103
use BUFX4  BUFX4_98
timestamp 1719641852
transform 1 0 1892 0 1 1905
box -2 -3 34 103
use OR2X2  OR2X2_20
timestamp 1719641852
transform 1 0 1924 0 1 1905
box -2 -3 34 103
use BUFX4  BUFX4_115
timestamp 1719641852
transform 1 0 1956 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_533
timestamp 1719641852
transform 1 0 1988 0 1 1905
box -2 -3 34 103
use DFFSR  DFFSR_184
timestamp 1719641852
transform -1 0 2196 0 1 1905
box -2 -3 178 103
use OAI21X1  OAI21X1_537
timestamp 1719641852
transform -1 0 2228 0 1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_184
timestamp 1719641852
transform -1 0 2260 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_534
timestamp 1719641852
transform -1 0 2292 0 1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_261
timestamp 1719641852
transform -1 0 2316 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_421
timestamp 1719641852
transform 1 0 2316 0 1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_137
timestamp 1719641852
transform 1 0 2348 0 1 1905
box -2 -3 34 103
use FILL  FILL_19_4_0
timestamp 1719641852
transform 1 0 2380 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_4_1
timestamp 1719641852
transform 1 0 2388 0 1 1905
box -2 -3 10 103
use AOI21X1  AOI21X1_117
timestamp 1719641852
transform 1 0 2396 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_369
timestamp 1719641852
transform -1 0 2460 0 1 1905
box -2 -3 34 103
use INVX2  INVX2_57
timestamp 1719641852
transform 1 0 2460 0 1 1905
box -2 -3 18 103
use OAI21X1  OAI21X1_470
timestamp 1719641852
transform -1 0 2508 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_469
timestamp 1719641852
transform -1 0 2540 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_425
timestamp 1719641852
transform -1 0 2572 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_317
timestamp 1719641852
transform 1 0 2572 0 1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_331
timestamp 1719641852
transform -1 0 2628 0 1 1905
box -2 -3 26 103
use AOI21X1  AOI21X1_255
timestamp 1719641852
transform -1 0 2660 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_762
timestamp 1719641852
transform -1 0 2692 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_761
timestamp 1719641852
transform -1 0 2724 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_760
timestamp 1719641852
transform 1 0 2724 0 1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_254
timestamp 1719641852
transform 1 0 2756 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_332
timestamp 1719641852
transform -1 0 2812 0 1 1905
box -2 -3 26 103
use BUFX4  BUFX4_135
timestamp 1719641852
transform 1 0 2812 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_778
timestamp 1719641852
transform 1 0 2844 0 1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_265
timestamp 1719641852
transform 1 0 2876 0 1 1905
box -2 -3 34 103
use FILL  FILL_19_5_0
timestamp 1719641852
transform -1 0 2916 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_5_1
timestamp 1719641852
transform -1 0 2924 0 1 1905
box -2 -3 10 103
use OAI21X1  OAI21X1_366
timestamp 1719641852
transform -1 0 2956 0 1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_113
timestamp 1719641852
transform -1 0 2988 0 1 1905
box -2 -3 34 103
use INVX2  INVX2_130
timestamp 1719641852
transform -1 0 3004 0 1 1905
box -2 -3 18 103
use NAND2X1  NAND2X1_225
timestamp 1719641852
transform 1 0 3004 0 1 1905
box -2 -3 26 103
use AOI22X1  AOI22X1_68
timestamp 1719641852
transform 1 0 3028 0 1 1905
box -2 -3 42 103
use OAI21X1  OAI21X1_307
timestamp 1719641852
transform 1 0 3068 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_305
timestamp 1719641852
transform 1 0 3100 0 1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_89
timestamp 1719641852
transform -1 0 3164 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_188
timestamp 1719641852
transform 1 0 3164 0 1 1905
box -2 -3 26 103
use AOI21X1  AOI21X1_91
timestamp 1719641852
transform -1 0 3220 0 1 1905
box -2 -3 34 103
use INVX1  INVX1_113
timestamp 1719641852
transform 1 0 3220 0 1 1905
box -2 -3 18 103
use NOR2X1  NOR2X1_189
timestamp 1719641852
transform -1 0 3260 0 1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_190
timestamp 1719641852
transform -1 0 3284 0 1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_146
timestamp 1719641852
transform 1 0 3284 0 1 1905
box -2 -3 26 103
use AOI21X1  AOI21X1_77
timestamp 1719641852
transform 1 0 3308 0 1 1905
box -2 -3 34 103
use AOI22X1  AOI22X1_51
timestamp 1719641852
transform 1 0 3340 0 1 1905
box -2 -3 42 103
use NAND2X1  NAND2X1_179
timestamp 1719641852
transform -1 0 3404 0 1 1905
box -2 -3 26 103
use FILL  FILL_19_6_0
timestamp 1719641852
transform -1 0 3412 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_6_1
timestamp 1719641852
transform -1 0 3420 0 1 1905
box -2 -3 10 103
use AOI21X1  AOI21X1_78
timestamp 1719641852
transform -1 0 3452 0 1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_147
timestamp 1719641852
transform 1 0 3452 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_250
timestamp 1719641852
transform 1 0 3476 0 1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_110
timestamp 1719641852
transform 1 0 3508 0 1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_109
timestamp 1719641852
transform 1 0 3532 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_225
timestamp 1719641852
transform 1 0 3556 0 1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_111
timestamp 1719641852
transform 1 0 3588 0 1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_112
timestamp 1719641852
transform 1 0 3612 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_226
timestamp 1719641852
transform -1 0 3668 0 1 1905
box -2 -3 34 103
use BUFX4  BUFX4_219
timestamp 1719641852
transform -1 0 3700 0 1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_166
timestamp 1719641852
transform -1 0 3732 0 1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_138
timestamp 1719641852
transform 1 0 3732 0 1 1905
box -2 -3 34 103
use FILL  FILL_20_1
timestamp 1719641852
transform 1 0 3764 0 1 1905
box -2 -3 10 103
use FILL  FILL_20_2
timestamp 1719641852
transform 1 0 3772 0 1 1905
box -2 -3 10 103
use BUFX2  BUFX2_16
timestamp 1719641852
transform -1 0 28 0 -1 2105
box -2 -3 26 103
use BUFX2  BUFX2_15
timestamp 1719641852
transform -1 0 52 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_139
timestamp 1719641852
transform 1 0 52 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_140
timestamp 1719641852
transform 1 0 84 0 -1 2105
box -2 -3 34 103
use DFFSR  DFFSR_14
timestamp 1719641852
transform -1 0 292 0 -1 2105
box -2 -3 178 103
use FILL  FILL_20_0_0
timestamp 1719641852
transform -1 0 300 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_0_1
timestamp 1719641852
transform -1 0 308 0 -1 2105
box -2 -3 10 103
use DFFSR  DFFSR_13
timestamp 1719641852
transform -1 0 484 0 -1 2105
box -2 -3 178 103
use INVX2  INVX2_5
timestamp 1719641852
transform 1 0 484 0 -1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_42
timestamp 1719641852
transform 1 0 500 0 -1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_40
timestamp 1719641852
transform 1 0 532 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_71
timestamp 1719641852
transform 1 0 564 0 -1 2105
box -2 -3 34 103
use INVX1  INVX1_20
timestamp 1719641852
transform 1 0 596 0 -1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_75
timestamp 1719641852
transform 1 0 612 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_33
timestamp 1719641852
transform -1 0 676 0 -1 2105
box -2 -3 34 103
use DFFSR  DFFSR_43
timestamp 1719641852
transform 1 0 676 0 -1 2105
box -2 -3 178 103
use FILL  FILL_20_1_0
timestamp 1719641852
transform 1 0 852 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_1_1
timestamp 1719641852
transform 1 0 860 0 -1 2105
box -2 -3 10 103
use OAI21X1  OAI21X1_68
timestamp 1719641852
transform 1 0 868 0 -1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_37
timestamp 1719641852
transform -1 0 932 0 -1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_85
timestamp 1719641852
transform -1 0 964 0 -1 2105
box -2 -3 34 103
use DFFSR  DFFSR_44
timestamp 1719641852
transform 1 0 964 0 -1 2105
box -2 -3 178 103
use NAND3X1  NAND3X1_67
timestamp 1719641852
transform 1 0 1140 0 -1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_68
timestamp 1719641852
transform 1 0 1172 0 -1 2105
box -2 -3 34 103
use INVX2  INVX2_17
timestamp 1719641852
transform -1 0 1220 0 -1 2105
box -2 -3 18 103
use NOR2X1  NOR2X1_4
timestamp 1719641852
transform 1 0 1220 0 -1 2105
box -2 -3 26 103
use NOR2X1  NOR2X1_3
timestamp 1719641852
transform 1 0 1244 0 -1 2105
box -2 -3 26 103
use BUFX4  BUFX4_128
timestamp 1719641852
transform -1 0 1300 0 -1 2105
box -2 -3 34 103
use CLKBUF1  CLKBUF1_13
timestamp 1719641852
transform -1 0 1372 0 -1 2105
box -2 -3 74 103
use FILL  FILL_20_2_0
timestamp 1719641852
transform 1 0 1372 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_2_1
timestamp 1719641852
transform 1 0 1380 0 -1 2105
box -2 -3 10 103
use BUFX4  BUFX4_208
timestamp 1719641852
transform 1 0 1388 0 -1 2105
box -2 -3 34 103
use INVX2  INVX2_92
timestamp 1719641852
transform 1 0 1420 0 -1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_637
timestamp 1719641852
transform 1 0 1436 0 -1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_235
timestamp 1719641852
transform -1 0 1500 0 -1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_236
timestamp 1719641852
transform 1 0 1500 0 -1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_291
timestamp 1719641852
transform 1 0 1532 0 -1 2105
box -2 -3 26 103
use DFFSR  DFFSR_136
timestamp 1719641852
transform 1 0 1556 0 -1 2105
box -2 -3 178 103
use OAI21X1  OAI21X1_678
timestamp 1719641852
transform 1 0 1732 0 -1 2105
box -2 -3 34 103
use INVX2  INVX2_90
timestamp 1719641852
transform 1 0 1764 0 -1 2105
box -2 -3 18 103
use NAND2X1  NAND2X1_295
timestamp 1719641852
transform 1 0 1780 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_674
timestamp 1719641852
transform -1 0 1836 0 -1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_339
timestamp 1719641852
transform 1 0 1836 0 -1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_264
timestamp 1719641852
transform -1 0 1892 0 -1 2105
box -2 -3 34 103
use FILL  FILL_20_3_0
timestamp 1719641852
transform -1 0 1900 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_3_1
timestamp 1719641852
transform -1 0 1908 0 -1 2105
box -2 -3 10 103
use OAI21X1  OAI21X1_774
timestamp 1719641852
transform -1 0 1940 0 -1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_335
timestamp 1719641852
transform 1 0 1940 0 -1 2105
box -2 -3 26 103
use DFFSR  DFFSR_185
timestamp 1719641852
transform -1 0 2140 0 -1 2105
box -2 -3 178 103
use INVX2  INVX2_95
timestamp 1719641852
transform -1 0 2156 0 -1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_535
timestamp 1719641852
transform 1 0 2156 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_536
timestamp 1719641852
transform 1 0 2188 0 -1 2105
box -2 -3 34 103
use INVX8  INVX8_21
timestamp 1719641852
transform 1 0 2220 0 -1 2105
box -2 -3 42 103
use AOI21X1  AOI21X1_139
timestamp 1719641852
transform 1 0 2260 0 -1 2105
box -2 -3 34 103
use INVX2  INVX2_93
timestamp 1719641852
transform -1 0 2308 0 -1 2105
box -2 -3 18 103
use NOR2X1  NOR2X1_227
timestamp 1719641852
transform 1 0 2308 0 -1 2105
box -2 -3 26 103
use INVX2  INVX2_132
timestamp 1719641852
transform 1 0 2332 0 -1 2105
box -2 -3 18 103
use NOR2X1  NOR2X1_336
timestamp 1719641852
transform 1 0 2348 0 -1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_267
timestamp 1719641852
transform -1 0 2404 0 -1 2105
box -2 -3 34 103
use FILL  FILL_20_4_0
timestamp 1719641852
transform 1 0 2404 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_4_1
timestamp 1719641852
transform 1 0 2412 0 -1 2105
box -2 -3 10 103
use OAI21X1  OAI21X1_771
timestamp 1719641852
transform 1 0 2420 0 -1 2105
box -2 -3 34 103
use BUFX4  BUFX4_37
timestamp 1719641852
transform 1 0 2452 0 -1 2105
box -2 -3 34 103
use BUFX4  BUFX4_169
timestamp 1719641852
transform 1 0 2484 0 -1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_262
timestamp 1719641852
transform -1 0 2540 0 -1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_185
timestamp 1719641852
transform 1 0 2540 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_539
timestamp 1719641852
transform 1 0 2572 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_764
timestamp 1719641852
transform 1 0 2604 0 -1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_256
timestamp 1719641852
transform -1 0 2668 0 -1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_51
timestamp 1719641852
transform -1 0 2692 0 -1 2105
box -2 -3 26 103
use AND2X2  AND2X2_32
timestamp 1719641852
transform -1 0 2724 0 -1 2105
box -2 -3 34 103
use INVX2  INVX2_77
timestamp 1719641852
transform 1 0 2724 0 -1 2105
box -2 -3 18 103
use DFFSR  DFFSR_183
timestamp 1719641852
transform 1 0 2740 0 -1 2105
box -2 -3 178 103
use FILL  FILL_20_5_0
timestamp 1719641852
transform 1 0 2916 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_5_1
timestamp 1719641852
transform 1 0 2924 0 -1 2105
box -2 -3 10 103
use INVX2  INVX2_116
timestamp 1719641852
transform 1 0 2932 0 -1 2105
box -2 -3 18 103
use NOR2X1  NOR2X1_211
timestamp 1719641852
transform -1 0 2972 0 -1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_111
timestamp 1719641852
transform 1 0 2972 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_357
timestamp 1719641852
transform -1 0 3036 0 -1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_216
timestamp 1719641852
transform 1 0 3036 0 -1 2105
box -2 -3 26 103
use BUFX4  BUFX4_66
timestamp 1719641852
transform -1 0 3092 0 -1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_93
timestamp 1719641852
transform -1 0 3124 0 -1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_60
timestamp 1719641852
transform 1 0 3124 0 -1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_99
timestamp 1719641852
transform 1 0 3156 0 -1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_61
timestamp 1719641852
transform 1 0 3188 0 -1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_148
timestamp 1719641852
transform 1 0 3220 0 -1 2105
box -2 -3 26 103
use NOR2X1  NOR2X1_129
timestamp 1719641852
transform 1 0 3244 0 -1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_163
timestamp 1719641852
transform -1 0 3292 0 -1 2105
box -2 -3 26 103
use NOR2X1  NOR2X1_170
timestamp 1719641852
transform 1 0 3292 0 -1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_178
timestamp 1719641852
transform 1 0 3316 0 -1 2105
box -2 -3 26 103
use NOR2X1  NOR2X1_171
timestamp 1719641852
transform 1 0 3340 0 -1 2105
box -2 -3 26 103
use NOR2X1  NOR2X1_149
timestamp 1719641852
transform 1 0 3364 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_251
timestamp 1719641852
transform 1 0 3388 0 -1 2105
box -2 -3 34 103
use FILL  FILL_20_6_0
timestamp 1719641852
transform 1 0 3420 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_6_1
timestamp 1719641852
transform 1 0 3428 0 -1 2105
box -2 -3 10 103
use OAI21X1  OAI21X1_263
timestamp 1719641852
transform 1 0 3436 0 -1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_172
timestamp 1719641852
transform 1 0 3468 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_264
timestamp 1719641852
transform 1 0 3492 0 -1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_164
timestamp 1719641852
transform -1 0 3556 0 -1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_159
timestamp 1719641852
transform -1 0 3588 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_111
timestamp 1719641852
transform -1 0 3612 0 -1 2105
box -2 -3 26 103
use NAND3X1  NAND3X1_165
timestamp 1719641852
transform -1 0 3644 0 -1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_71
timestamp 1719641852
transform 1 0 3644 0 -1 2105
box -2 -3 26 103
use NAND3X1  NAND3X1_169
timestamp 1719641852
transform 1 0 3668 0 -1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_167
timestamp 1719641852
transform -1 0 3732 0 -1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_168
timestamp 1719641852
transform 1 0 3732 0 -1 2105
box -2 -3 34 103
use INVX1  INVX1_82
timestamp 1719641852
transform 1 0 3764 0 -1 2105
box -2 -3 18 103
use BUFX2  BUFX2_12
timestamp 1719641852
transform -1 0 28 0 1 2105
box -2 -3 26 103
use DFFSR  DFFSR_74
timestamp 1719641852
transform -1 0 204 0 1 2105
box -2 -3 178 103
use CLKBUF1  CLKBUF1_23
timestamp 1719641852
transform 1 0 204 0 1 2105
box -2 -3 74 103
use FILL  FILL_21_0_0
timestamp 1719641852
transform 1 0 276 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_0_1
timestamp 1719641852
transform 1 0 284 0 1 2105
box -2 -3 10 103
use DFFSR  DFFSR_45
timestamp 1719641852
transform 1 0 292 0 1 2105
box -2 -3 178 103
use BUFX4  BUFX4_140
timestamp 1719641852
transform -1 0 500 0 1 2105
box -2 -3 34 103
use INVX1  INVX1_19
timestamp 1719641852
transform 1 0 500 0 1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_72
timestamp 1719641852
transform 1 0 516 0 1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_39
timestamp 1719641852
transform -1 0 580 0 1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_19
timestamp 1719641852
transform 1 0 580 0 1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_25
timestamp 1719641852
transform 1 0 612 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_183
timestamp 1719641852
transform -1 0 676 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_182
timestamp 1719641852
transform 1 0 676 0 1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_36
timestamp 1719641852
transform -1 0 740 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_66
timestamp 1719641852
transform -1 0 772 0 1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_38
timestamp 1719641852
transform -1 0 804 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_70
timestamp 1719641852
transform -1 0 836 0 1 2105
box -2 -3 34 103
use FILL  FILL_21_1_0
timestamp 1719641852
transform -1 0 844 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_1_1
timestamp 1719641852
transform -1 0 852 0 1 2105
box -2 -3 10 103
use DFFSR  DFFSR_155
timestamp 1719641852
transform -1 0 1028 0 1 2105
box -2 -3 178 103
use CLKBUF1  CLKBUF1_5
timestamp 1719641852
transform 1 0 1028 0 1 2105
box -2 -3 74 103
use OAI21X1  OAI21X1_718
timestamp 1719641852
transform 1 0 1100 0 1 2105
box -2 -3 34 103
use INVX1  INVX1_43
timestamp 1719641852
transform -1 0 1148 0 1 2105
box -2 -3 18 103
use NAND2X1  NAND2X1_318
timestamp 1719641852
transform -1 0 1172 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_721
timestamp 1719641852
transform -1 0 1204 0 1 2105
box -2 -3 34 103
use DFFSR  DFFSR_152
timestamp 1719641852
transform -1 0 1380 0 1 2105
box -2 -3 178 103
use FILL  FILL_21_2_0
timestamp 1719641852
transform -1 0 1388 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_2_1
timestamp 1719641852
transform -1 0 1396 0 1 2105
box -2 -3 10 103
use INVX1  INVX1_36
timestamp 1719641852
transform -1 0 1412 0 1 2105
box -2 -3 18 103
use INVX8  INVX8_22
timestamp 1719641852
transform -1 0 1452 0 1 2105
box -2 -3 42 103
use AOI22X1  AOI22X1_8
timestamp 1719641852
transform 1 0 1452 0 1 2105
box -2 -3 42 103
use NAND2X1  NAND2X1_338
timestamp 1719641852
transform 1 0 1492 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_784
timestamp 1719641852
transform 1 0 1516 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_783
timestamp 1719641852
transform -1 0 1580 0 1 2105
box -2 -3 34 103
use INVX1  INVX1_164
timestamp 1719641852
transform 1 0 1580 0 1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_788
timestamp 1719641852
transform 1 0 1596 0 1 2105
box -2 -3 34 103
use INVX2  INVX2_133
timestamp 1719641852
transform 1 0 1628 0 1 2105
box -2 -3 18 103
use NAND2X1  NAND2X1_336
timestamp 1719641852
transform 1 0 1644 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_777
timestamp 1719641852
transform -1 0 1700 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_776
timestamp 1719641852
transform -1 0 1732 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_775
timestamp 1719641852
transform -1 0 1764 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_33
timestamp 1719641852
transform -1 0 1796 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_528
timestamp 1719641852
transform 1 0 1796 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_532
timestamp 1719641852
transform -1 0 1860 0 1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_183
timestamp 1719641852
transform -1 0 1892 0 1 2105
box -2 -3 34 103
use FILL  FILL_21_3_0
timestamp 1719641852
transform 1 0 1892 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_3_1
timestamp 1719641852
transform 1 0 1900 0 1 2105
box -2 -3 10 103
use OAI21X1  OAI21X1_529
timestamp 1719641852
transform 1 0 1908 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_531
timestamp 1719641852
transform 1 0 1940 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_530
timestamp 1719641852
transform -1 0 2004 0 1 2105
box -2 -3 34 103
use DFFSR  DFFSR_219
timestamp 1719641852
transform -1 0 2180 0 1 2105
box -2 -3 178 103
use AND2X2  AND2X2_26
timestamp 1719641852
transform -1 0 2212 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_422
timestamp 1719641852
transform -1 0 2244 0 1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_138
timestamp 1719641852
transform 1 0 2244 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_779
timestamp 1719641852
transform -1 0 2308 0 1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_266
timestamp 1719641852
transform 1 0 2308 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_413
timestamp 1719641852
transform -1 0 2372 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_540
timestamp 1719641852
transform -1 0 2404 0 1 2105
box -2 -3 34 103
use FILL  FILL_21_4_0
timestamp 1719641852
transform 1 0 2404 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_4_1
timestamp 1719641852
transform 1 0 2412 0 1 2105
box -2 -3 10 103
use OAI21X1  OAI21X1_541
timestamp 1719641852
transform 1 0 2420 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_538
timestamp 1719641852
transform 1 0 2452 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_763
timestamp 1719641852
transform 1 0 2484 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_542
timestamp 1719641852
transform -1 0 2548 0 1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_249
timestamp 1719641852
transform 1 0 2548 0 1 2105
box -2 -3 26 103
use BUFX4  BUFX4_48
timestamp 1719641852
transform -1 0 2604 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_47
timestamp 1719641852
transform 1 0 2604 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_418
timestamp 1719641852
transform -1 0 2668 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_372
timestamp 1719641852
transform -1 0 2700 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_358
timestamp 1719641852
transform -1 0 2732 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_359
timestamp 1719641852
transform 1 0 2732 0 1 2105
box -2 -3 34 103
use INVX2  INVX2_52
timestamp 1719641852
transform -1 0 2780 0 1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_356
timestamp 1719641852
transform 1 0 2780 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_360
timestamp 1719641852
transform -1 0 2844 0 1 2105
box -2 -3 34 103
use FILL  FILL_21_5_0
timestamp 1719641852
transform -1 0 2852 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_5_1
timestamp 1719641852
transform -1 0 2860 0 1 2105
box -2 -3 10 103
use DFFSR  DFFSR_234
timestamp 1719641852
transform -1 0 3036 0 1 2105
box -2 -3 178 103
use OR2X2  OR2X2_13
timestamp 1719641852
transform -1 0 3068 0 1 2105
box -2 -3 34 103
use OR2X2  OR2X2_12
timestamp 1719641852
transform -1 0 3100 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_161
timestamp 1719641852
transform 1 0 3100 0 1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_98
timestamp 1719641852
transform 1 0 3124 0 1 2105
box -2 -3 34 103
use AOI22X1  AOI22X1_42
timestamp 1719641852
transform 1 0 3156 0 1 2105
box -2 -3 42 103
use OAI21X1  OAI21X1_296
timestamp 1719641852
transform -1 0 3228 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_164
timestamp 1719641852
transform 1 0 3228 0 1 2105
box -2 -3 26 103
use AOI22X1  AOI22X1_43
timestamp 1719641852
transform 1 0 3252 0 1 2105
box -2 -3 42 103
use NAND2X1  NAND2X1_162
timestamp 1719641852
transform -1 0 3316 0 1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_94
timestamp 1719641852
transform -1 0 3348 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_157
timestamp 1719641852
transform -1 0 3380 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_178
timestamp 1719641852
transform -1 0 3412 0 1 2105
box -2 -3 34 103
use FILL  FILL_21_6_0
timestamp 1719641852
transform 1 0 3412 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_6_1
timestamp 1719641852
transform 1 0 3420 0 1 2105
box -2 -3 10 103
use NOR2X1  NOR2X1_173
timestamp 1719641852
transform 1 0 3428 0 1 2105
box -2 -3 26 103
use NOR2X1  NOR2X1_169
timestamp 1719641852
transform -1 0 3476 0 1 2105
box -2 -3 26 103
use NOR2X1  NOR2X1_168
timestamp 1719641852
transform 1 0 3476 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_262
timestamp 1719641852
transform 1 0 3500 0 1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_95
timestamp 1719641852
transform 1 0 3532 0 1 2105
box -2 -3 26 103
use NAND3X1  NAND3X1_110
timestamp 1719641852
transform -1 0 3588 0 1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_109
timestamp 1719641852
transform -1 0 3620 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_42
timestamp 1719641852
transform -1 0 3652 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_213
timestamp 1719641852
transform -1 0 3684 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_206
timestamp 1719641852
transform 1 0 3684 0 1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_112
timestamp 1719641852
transform 1 0 3716 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_185
timestamp 1719641852
transform -1 0 3780 0 1 2105
box -2 -3 34 103
use BUFX2  BUFX2_11
timestamp 1719641852
transform -1 0 28 0 -1 2305
box -2 -3 26 103
use CLKBUF1  CLKBUF1_55
timestamp 1719641852
transform 1 0 28 0 -1 2305
box -2 -3 74 103
use OAI21X1  OAI21X1_135
timestamp 1719641852
transform 1 0 100 0 -1 2305
box -2 -3 34 103
use CLKBUF1  CLKBUF1_40
timestamp 1719641852
transform 1 0 132 0 -1 2305
box -2 -3 74 103
use BUFX4  BUFX4_102
timestamp 1719641852
transform -1 0 236 0 -1 2305
box -2 -3 34 103
use DFFSR  DFFSR_9
timestamp 1719641852
transform -1 0 412 0 -1 2305
box -2 -3 178 103
use FILL  FILL_22_0_0
timestamp 1719641852
transform 1 0 412 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_0_1
timestamp 1719641852
transform 1 0 420 0 -1 2305
box -2 -3 10 103
use INVX2  INVX2_1
timestamp 1719641852
transform 1 0 428 0 -1 2305
box -2 -3 18 103
use OAI21X1  OAI21X1_34
timestamp 1719641852
transform 1 0 444 0 -1 2305
box -2 -3 34 103
use DFFSR  DFFSR_47
timestamp 1719641852
transform -1 0 652 0 -1 2305
box -2 -3 178 103
use DFFSR  DFFSR_53
timestamp 1719641852
transform -1 0 828 0 -1 2305
box -2 -3 178 103
use BUFX4  BUFX4_27
timestamp 1719641852
transform -1 0 860 0 -1 2305
box -2 -3 34 103
use FILL  FILL_22_1_0
timestamp 1719641852
transform -1 0 868 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_1_1
timestamp 1719641852
transform -1 0 876 0 -1 2305
box -2 -3 10 103
use BUFX4  BUFX4_18
timestamp 1719641852
transform -1 0 908 0 -1 2305
box -2 -3 34 103
use BUFX4  BUFX4_201
timestamp 1719641852
transform 1 0 908 0 -1 2305
box -2 -3 34 103
use OAI22X1  OAI22X1_20
timestamp 1719641852
transform 1 0 940 0 -1 2305
box -2 -3 42 103
use INVX1  INVX1_45
timestamp 1719641852
transform -1 0 996 0 -1 2305
box -2 -3 18 103
use NOR2X1  NOR2X1_11
timestamp 1719641852
transform -1 0 1020 0 -1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_47
timestamp 1719641852
transform -1 0 1044 0 -1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_8
timestamp 1719641852
transform -1 0 1076 0 -1 2305
box -2 -3 34 103
use OAI22X1  OAI22X1_19
timestamp 1719641852
transform 1 0 1076 0 -1 2305
box -2 -3 42 103
use INVX2  INVX2_94
timestamp 1719641852
transform 1 0 1116 0 -1 2305
box -2 -3 18 103
use BUFX4  BUFX4_225
timestamp 1719641852
transform 1 0 1132 0 -1 2305
box -2 -3 34 103
use INVX1  INVX1_44
timestamp 1719641852
transform -1 0 1180 0 -1 2305
box -2 -3 18 103
use NAND3X1  NAND3X1_76
timestamp 1719641852
transform 1 0 1180 0 -1 2305
box -2 -3 34 103
use DFFSR  DFFSR_122
timestamp 1719641852
transform -1 0 1388 0 -1 2305
box -2 -3 178 103
use FILL  FILL_22_2_0
timestamp 1719641852
transform 1 0 1388 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_2_1
timestamp 1719641852
transform 1 0 1396 0 -1 2305
box -2 -3 10 103
use INVX2  INVX2_60
timestamp 1719641852
transform 1 0 1404 0 -1 2305
box -2 -3 18 103
use OAI21X1  OAI21X1_714
timestamp 1719641852
transform -1 0 1452 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_315
timestamp 1719641852
transform 1 0 1452 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_713
timestamp 1719641852
transform -1 0 1508 0 -1 2305
box -2 -3 34 103
use INVX2  INVX2_135
timestamp 1719641852
transform 1 0 1508 0 -1 2305
box -2 -3 18 103
use DFFSR  DFFSR_123
timestamp 1719641852
transform -1 0 1700 0 -1 2305
box -2 -3 178 103
use OAI21X1  OAI21X1_789
timestamp 1719641852
transform -1 0 1732 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_341
timestamp 1719641852
transform -1 0 1756 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_711
timestamp 1719641852
transform -1 0 1788 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_712
timestamp 1719641852
transform -1 0 1820 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_314
timestamp 1719641852
transform -1 0 1844 0 -1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_290
timestamp 1719641852
transform -1 0 1868 0 -1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_289
timestamp 1719641852
transform 1 0 1868 0 -1 2305
box -2 -3 26 103
use FILL  FILL_22_3_0
timestamp 1719641852
transform 1 0 1892 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_3_1
timestamp 1719641852
transform 1 0 1900 0 -1 2305
box -2 -3 10 103
use INVX2  INVX2_58
timestamp 1719641852
transform 1 0 1908 0 -1 2305
box -2 -3 18 103
use AOI21X1  AOI21X1_230
timestamp 1719641852
transform -1 0 1956 0 -1 2305
box -2 -3 34 103
use INVX2  INVX2_157
timestamp 1719641852
transform 1 0 1956 0 -1 2305
box -2 -3 18 103
use AOI21X1  AOI21X1_231
timestamp 1719641852
transform -1 0 2004 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_631
timestamp 1719641852
transform -1 0 2036 0 -1 2305
box -2 -3 34 103
use BUFX4  BUFX4_28
timestamp 1719641852
transform -1 0 2068 0 -1 2305
box -2 -3 34 103
use BUFX4  BUFX4_32
timestamp 1719641852
transform 1 0 2068 0 -1 2305
box -2 -3 34 103
use BUFX4  BUFX4_60
timestamp 1719641852
transform 1 0 2100 0 -1 2305
box -2 -3 34 103
use INVX8  INVX8_20
timestamp 1719641852
transform 1 0 2132 0 -1 2305
box -2 -3 42 103
use DFFSR  DFFSR_216
timestamp 1719641852
transform -1 0 2348 0 -1 2305
box -2 -3 178 103
use OAI21X1  OAI21X1_525
timestamp 1719641852
transform -1 0 2380 0 -1 2305
box -2 -3 34 103
use FILL  FILL_22_4_0
timestamp 1719641852
transform -1 0 2388 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_4_1
timestamp 1719641852
transform -1 0 2396 0 -1 2305
box -2 -3 10 103
use OAI21X1  OAI21X1_526
timestamp 1719641852
transform -1 0 2428 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_765
timestamp 1719641852
transform -1 0 2460 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_766
timestamp 1719641852
transform 1 0 2460 0 -1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_182
timestamp 1719641852
transform 1 0 2492 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_524
timestamp 1719641852
transform -1 0 2556 0 -1 2305
box -2 -3 34 103
use AND2X2  AND2X2_25
timestamp 1719641852
transform -1 0 2588 0 -1 2305
box -2 -3 34 103
use AND2X2  AND2X2_27
timestamp 1719641852
transform -1 0 2620 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_767
timestamp 1719641852
transform -1 0 2652 0 -1 2305
box -2 -3 34 103
use DFFSR  DFFSR_187
timestamp 1719641852
transform 1 0 2652 0 -1 2305
box -2 -3 178 103
use NOR2X1  NOR2X1_243
timestamp 1719641852
transform 1 0 2828 0 -1 2305
box -2 -3 26 103
use BUFX4  BUFX4_151
timestamp 1719641852
transform -1 0 2884 0 -1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_253
timestamp 1719641852
transform 1 0 2884 0 -1 2305
box -2 -3 26 103
use FILL  FILL_22_5_0
timestamp 1719641852
transform -1 0 2916 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_5_1
timestamp 1719641852
transform -1 0 2924 0 -1 2305
box -2 -3 10 103
use INVX2  INVX2_134
timestamp 1719641852
transform -1 0 2940 0 -1 2305
box -2 -3 18 103
use BUFX4  BUFX4_152
timestamp 1719641852
transform -1 0 2972 0 -1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_144
timestamp 1719641852
transform -1 0 3004 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_430
timestamp 1719641852
transform -1 0 3036 0 -1 2305
box -2 -3 34 103
use INVX2  INVX2_59
timestamp 1719641852
transform 1 0 3036 0 -1 2305
box -2 -3 18 103
use AOI21X1  AOI21X1_101
timestamp 1719641852
transform 1 0 3052 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_313
timestamp 1719641852
transform -1 0 3116 0 -1 2305
box -2 -3 34 103
use NAND3X1  NAND3X1_208
timestamp 1719641852
transform 1 0 3116 0 -1 2305
box -2 -3 34 103
use AOI22X1  AOI22X1_67
timestamp 1719641852
transform 1 0 3148 0 -1 2305
box -2 -3 42 103
use NAND2X1  NAND2X1_196
timestamp 1719641852
transform -1 0 3212 0 -1 2305
box -2 -3 26 103
use AOI22X1  AOI22X1_66
timestamp 1719641852
transform -1 0 3252 0 -1 2305
box -2 -3 42 103
use NAND2X1  NAND2X1_193
timestamp 1719641852
transform -1 0 3276 0 -1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_62
timestamp 1719641852
transform -1 0 3308 0 -1 2305
box -2 -3 34 103
use BUFX4  BUFX4_176
timestamp 1719641852
transform -1 0 3340 0 -1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_70
timestamp 1719641852
transform 1 0 3340 0 -1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_69
timestamp 1719641852
transform 1 0 3364 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_205
timestamp 1719641852
transform 1 0 3388 0 -1 2305
box -2 -3 34 103
use FILL  FILL_22_6_0
timestamp 1719641852
transform 1 0 3420 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_6_1
timestamp 1719641852
transform 1 0 3428 0 -1 2305
box -2 -3 10 103
use NOR2X1  NOR2X1_73
timestamp 1719641852
transform 1 0 3436 0 -1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_74
timestamp 1719641852
transform 1 0 3460 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_207
timestamp 1719641852
transform 1 0 3484 0 -1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_96
timestamp 1719641852
transform 1 0 3516 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_218
timestamp 1719641852
transform 1 0 3540 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_113
timestamp 1719641852
transform 1 0 3572 0 -1 2305
box -2 -3 26 103
use NAND3X1  NAND3X1_163
timestamp 1719641852
transform -1 0 3628 0 -1 2305
box -2 -3 34 103
use NAND3X1  NAND3X1_121
timestamp 1719641852
transform -1 0 3660 0 -1 2305
box -2 -3 34 103
use NAND3X1  NAND3X1_122
timestamp 1719641852
transform -1 0 3692 0 -1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_72
timestamp 1719641852
transform 1 0 3692 0 -1 2305
box -2 -3 26 103
use NAND3X1  NAND3X1_111
timestamp 1719641852
transform -1 0 3748 0 -1 2305
box -2 -3 34 103
use BUFX4  BUFX4_239
timestamp 1719641852
transform -1 0 3780 0 -1 2305
box -2 -3 34 103
use BUFX2  BUFX2_45
timestamp 1719641852
transform -1 0 28 0 1 2305
box -2 -3 26 103
use BUFX2  BUFX2_43
timestamp 1719641852
transform -1 0 52 0 1 2305
box -2 -3 26 103
use DFFSR  DFFSR_72
timestamp 1719641852
transform -1 0 228 0 1 2305
box -2 -3 178 103
use DFFSR  DFFSR_54
timestamp 1719641852
transform 1 0 228 0 1 2305
box -2 -3 178 103
use FILL  FILL_23_0_0
timestamp 1719641852
transform 1 0 404 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_0_1
timestamp 1719641852
transform 1 0 412 0 1 2305
box -2 -3 10 103
use INVX2  INVX2_38
timestamp 1719641852
transform 1 0 420 0 1 2305
box -2 -3 18 103
use INVX2  INVX2_7
timestamp 1719641852
transform 1 0 436 0 1 2305
box -2 -3 18 103
use BUFX4  BUFX4_142
timestamp 1719641852
transform 1 0 452 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_46
timestamp 1719641852
transform 1 0 484 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_125
timestamp 1719641852
transform 1 0 516 0 1 2305
box -2 -3 34 103
use INVX2  INVX2_31
timestamp 1719641852
transform 1 0 548 0 1 2305
box -2 -3 18 103
use OAI21X1  OAI21X1_111
timestamp 1719641852
transform 1 0 564 0 1 2305
box -2 -3 34 103
use NAND3X1  NAND3X1_66
timestamp 1719641852
transform 1 0 596 0 1 2305
box -2 -3 34 103
use BUFX4  BUFX4_106
timestamp 1719641852
transform -1 0 660 0 1 2305
box -2 -3 34 103
use INVX2  INVX2_37
timestamp 1719641852
transform 1 0 660 0 1 2305
box -2 -3 18 103
use OAI21X1  OAI21X1_124
timestamp 1719641852
transform 1 0 676 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_123
timestamp 1719641852
transform 1 0 708 0 1 2305
box -2 -3 34 103
use NAND3X1  NAND3X1_65
timestamp 1719641852
transform 1 0 740 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_333
timestamp 1719641852
transform 1 0 772 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_122
timestamp 1719641852
transform 1 0 796 0 1 2305
box -2 -3 34 103
use INVX8  INVX8_1
timestamp 1719641852
transform -1 0 868 0 1 2305
box -2 -3 42 103
use FILL  FILL_23_1_0
timestamp 1719641852
transform -1 0 876 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_1_1
timestamp 1719641852
transform -1 0 884 0 1 2305
box -2 -3 10 103
use OAI22X1  OAI22X1_16
timestamp 1719641852
transform -1 0 924 0 1 2305
box -2 -3 42 103
use INVX1  INVX1_28
timestamp 1719641852
transform -1 0 940 0 1 2305
box -2 -3 18 103
use BUFX4  BUFX4_75
timestamp 1719641852
transform -1 0 972 0 1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_10
timestamp 1719641852
transform 1 0 972 0 1 2305
box -2 -3 26 103
use BUFX4  BUFX4_228
timestamp 1719641852
transform -1 0 1028 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_46
timestamp 1719641852
transform -1 0 1052 0 1 2305
box -2 -3 26 103
use DFFSR  DFFSR_120
timestamp 1719641852
transform -1 0 1228 0 1 2305
box -2 -3 178 103
use INVX1  INVX1_35
timestamp 1719641852
transform 1 0 1228 0 1 2305
box -2 -3 18 103
use OAI22X1  OAI22X1_11
timestamp 1719641852
transform 1 0 1244 0 1 2305
box -2 -3 42 103
use OAI22X1  OAI22X1_17
timestamp 1719641852
transform 1 0 1284 0 1 2305
box -2 -3 42 103
use INVX1  INVX1_41
timestamp 1719641852
transform -1 0 1340 0 1 2305
box -2 -3 18 103
use INVX1  INVX1_42
timestamp 1719641852
transform -1 0 1356 0 1 2305
box -2 -3 18 103
use FILL  FILL_23_2_0
timestamp 1719641852
transform -1 0 1364 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_2_1
timestamp 1719641852
transform -1 0 1372 0 1 2305
box -2 -3 10 103
use DFFSR  DFFSR_154
timestamp 1719641852
transform -1 0 1548 0 1 2305
box -2 -3 178 103
use OAI21X1  OAI21X1_786
timestamp 1719641852
transform 1 0 1548 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_787
timestamp 1719641852
transform 1 0 1580 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_340
timestamp 1719641852
transform -1 0 1636 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_790
timestamp 1719641852
transform -1 0 1668 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_339
timestamp 1719641852
transform -1 0 1692 0 1 2305
box -2 -3 26 103
use BUFX4  BUFX4_206
timestamp 1719641852
transform 1 0 1692 0 1 2305
box -2 -3 34 103
use INVX1  INVX1_37
timestamp 1719641852
transform -1 0 1740 0 1 2305
box -2 -3 18 103
use INVX1  INVX1_39
timestamp 1719641852
transform -1 0 1756 0 1 2305
box -2 -3 18 103
use INVX1  INVX1_33
timestamp 1719641852
transform -1 0 1772 0 1 2305
box -2 -3 18 103
use OAI21X1  OAI21X1_667
timestamp 1719641852
transform 1 0 1772 0 1 2305
box -2 -3 34 103
use INVX1  INVX1_149
timestamp 1719641852
transform -1 0 1820 0 1 2305
box -2 -3 18 103
use OAI21X1  OAI21X1_668
timestamp 1719641852
transform -1 0 1852 0 1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_307
timestamp 1719641852
transform 1 0 1852 0 1 2305
box -2 -3 26 103
use FILL  FILL_23_3_0
timestamp 1719641852
transform -1 0 1884 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_3_1
timestamp 1719641852
transform -1 0 1892 0 1 2305
box -2 -3 10 103
use AOI21X1  AOI21X1_232
timestamp 1719641852
transform -1 0 1924 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_630
timestamp 1719641852
transform -1 0 1956 0 1 2305
box -2 -3 34 103
use OR2X2  OR2X2_17
timestamp 1719641852
transform -1 0 1988 0 1 2305
box -2 -3 34 103
use INVX1  INVX1_34
timestamp 1719641852
transform -1 0 2004 0 1 2305
box -2 -3 18 103
use OAI21X1  OAI21X1_523
timestamp 1719641852
transform 1 0 2004 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_585
timestamp 1719641852
transform 1 0 2036 0 1 2305
box -2 -3 34 103
use DFFSR  DFFSR_212
timestamp 1719641852
transform -1 0 2244 0 1 2305
box -2 -3 178 103
use BUFX4  BUFX4_171
timestamp 1719641852
transform 1 0 2244 0 1 2305
box -2 -3 34 103
use BUFX4  BUFX4_170
timestamp 1719641852
transform 1 0 2276 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_527
timestamp 1719641852
transform -1 0 2340 0 1 2305
box -2 -3 34 103
use FILL  FILL_23_4_0
timestamp 1719641852
transform 1 0 2340 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_4_1
timestamp 1719641852
transform 1 0 2348 0 1 2305
box -2 -3 10 103
use DFFSR  DFFSR_186
timestamp 1719641852
transform 1 0 2356 0 1 2305
box -2 -3 178 103
use OAI21X1  OAI21X1_433
timestamp 1719641852
transform -1 0 2564 0 1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_231
timestamp 1719641852
transform 1 0 2564 0 1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_149
timestamp 1719641852
transform -1 0 2620 0 1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_148
timestamp 1719641852
transform -1 0 2652 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_432
timestamp 1719641852
transform 1 0 2652 0 1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_147
timestamp 1719641852
transform 1 0 2684 0 1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_251
timestamp 1719641852
transform 1 0 2716 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_380
timestamp 1719641852
transform 1 0 2740 0 1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_121
timestamp 1719641852
transform -1 0 2804 0 1 2305
box -2 -3 34 103
use INVX2  INVX2_145
timestamp 1719641852
transform 1 0 2804 0 1 2305
box -2 -3 18 103
use NOR2X1  NOR2X1_230
timestamp 1719641852
transform 1 0 2820 0 1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_146
timestamp 1719641852
transform -1 0 2876 0 1 2305
box -2 -3 34 103
use FILL  FILL_23_5_0
timestamp 1719641852
transform -1 0 2884 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_5_1
timestamp 1719641852
transform -1 0 2892 0 1 2305
box -2 -3 10 103
use DFFSR  DFFSR_213
timestamp 1719641852
transform -1 0 3068 0 1 2305
box -2 -3 178 103
use AOI21X1  AOI21X1_100
timestamp 1719641852
transform 1 0 3068 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_312
timestamp 1719641852
transform -1 0 3132 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_195
timestamp 1719641852
transform 1 0 3132 0 1 2305
box -2 -3 26 103
use INVX1  INVX1_117
timestamp 1719641852
transform 1 0 3156 0 1 2305
box -2 -3 18 103
use AOI22X1  AOI22X1_37
timestamp 1719641852
transform 1 0 3172 0 1 2305
box -2 -3 42 103
use NAND2X1  NAND2X1_155
timestamp 1719641852
transform 1 0 3212 0 1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_52
timestamp 1719641852
transform -1 0 3268 0 1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_95
timestamp 1719641852
transform -1 0 3300 0 1 2305
box -2 -3 34 103
use BUFX4  BUFX4_154
timestamp 1719641852
transform -1 0 3332 0 1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_98
timestamp 1719641852
transform 1 0 3332 0 1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_97
timestamp 1719641852
transform 1 0 3356 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_219
timestamp 1719641852
transform 1 0 3380 0 1 2305
box -2 -3 34 103
use FILL  FILL_23_6_0
timestamp 1719641852
transform -1 0 3420 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_6_1
timestamp 1719641852
transform -1 0 3428 0 1 2305
box -2 -3 10 103
use NAND3X1  NAND3X1_157
timestamp 1719641852
transform -1 0 3460 0 1 2305
box -2 -3 34 103
use NAND3X1  NAND3X1_158
timestamp 1719641852
transform 1 0 3460 0 1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_166
timestamp 1719641852
transform 1 0 3492 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_261
timestamp 1719641852
transform 1 0 3516 0 1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_115
timestamp 1719641852
transform 1 0 3548 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_234
timestamp 1719641852
transform 1 0 3572 0 1 2305
box -2 -3 34 103
use NAND3X1  NAND3X1_136
timestamp 1719641852
transform -1 0 3636 0 1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_113
timestamp 1719641852
transform 1 0 3636 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_233
timestamp 1719641852
transform 1 0 3660 0 1 2305
box -2 -3 34 103
use NAND3X1  NAND3X1_135
timestamp 1719641852
transform -1 0 3724 0 1 2305
box -2 -3 34 103
use NAND3X1  NAND3X1_137
timestamp 1719641852
transform -1 0 3756 0 1 2305
box -2 -3 34 103
use FILL  FILL_24_1
timestamp 1719641852
transform 1 0 3756 0 1 2305
box -2 -3 10 103
use FILL  FILL_24_2
timestamp 1719641852
transform 1 0 3764 0 1 2305
box -2 -3 10 103
use FILL  FILL_24_3
timestamp 1719641852
transform 1 0 3772 0 1 2305
box -2 -3 10 103
use BUFX2  BUFX2_55
timestamp 1719641852
transform -1 0 28 0 -1 2505
box -2 -3 26 103
use BUFX2  BUFX2_10
timestamp 1719641852
transform -1 0 52 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_134
timestamp 1719641852
transform 1 0 52 0 -1 2505
box -2 -3 34 103
use DFFSR  DFFSR_84
timestamp 1719641852
transform -1 0 260 0 -1 2505
box -2 -3 178 103
use FILL  FILL_24_0_0
timestamp 1719641852
transform -1 0 268 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_0_1
timestamp 1719641852
transform -1 0 276 0 -1 2505
box -2 -3 10 103
use DFFSR  DFFSR_8
timestamp 1719641852
transform -1 0 452 0 -1 2505
box -2 -3 178 103
use INVX2  INVX2_16
timestamp 1719641852
transform 1 0 452 0 -1 2505
box -2 -3 18 103
use DFFSR  DFFSR_50
timestamp 1719641852
transform 1 0 468 0 -1 2505
box -2 -3 178 103
use NAND3X1  NAND3X1_59
timestamp 1719641852
transform 1 0 644 0 -1 2505
box -2 -3 34 103
use INVX2  INVX2_34
timestamp 1719641852
transform 1 0 676 0 -1 2505
box -2 -3 18 103
use BUFX4  BUFX4_107
timestamp 1719641852
transform 1 0 692 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_117
timestamp 1719641852
transform 1 0 724 0 -1 2505
box -2 -3 34 103
use NAND3X1  NAND3X1_62
timestamp 1719641852
transform -1 0 788 0 -1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_32
timestamp 1719641852
transform -1 0 812 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_116
timestamp 1719641852
transform -1 0 844 0 -1 2505
box -2 -3 34 103
use FILL  FILL_24_1_0
timestamp 1719641852
transform -1 0 852 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_1_1
timestamp 1719641852
transform -1 0 860 0 -1 2505
box -2 -3 10 103
use BUFX4  BUFX4_13
timestamp 1719641852
transform -1 0 892 0 -1 2505
box -2 -3 34 103
use OAI22X1  OAI22X1_7
timestamp 1719641852
transform -1 0 932 0 -1 2505
box -2 -3 42 103
use OAI22X1  OAI22X1_10
timestamp 1719641852
transform -1 0 972 0 -1 2505
box -2 -3 42 103
use NAND2X1  NAND2X1_45
timestamp 1719641852
transform -1 0 996 0 -1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_8
timestamp 1719641852
transform 1 0 996 0 -1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_43
timestamp 1719641852
transform -1 0 1044 0 -1 2505
box -2 -3 26 103
use BUFX4  BUFX4_78
timestamp 1719641852
transform 1 0 1044 0 -1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_5
timestamp 1719641852
transform 1 0 1076 0 -1 2505
box -2 -3 34 103
use OAI22X1  OAI22X1_12
timestamp 1719641852
transform -1 0 1148 0 -1 2505
box -2 -3 42 103
use AOI21X1  AOI21X1_7
timestamp 1719641852
transform -1 0 1180 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_7
timestamp 1719641852
transform 1 0 1180 0 -1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_127
timestamp 1719641852
transform 1 0 1204 0 -1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_42
timestamp 1719641852
transform -1 0 1252 0 -1 2505
box -2 -3 26 103
use AOI21X1  AOI21X1_4
timestamp 1719641852
transform -1 0 1284 0 -1 2505
box -2 -3 34 103
use CLKBUF1  CLKBUF1_51
timestamp 1719641852
transform 1 0 1284 0 -1 2505
box -2 -3 74 103
use FILL  FILL_24_2_0
timestamp 1719641852
transform -1 0 1364 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_2_1
timestamp 1719641852
transform -1 0 1372 0 -1 2505
box -2 -3 10 103
use INVX8  INVX8_5
timestamp 1719641852
transform -1 0 1412 0 -1 2505
box -2 -3 42 103
use BUFX4  BUFX4_191
timestamp 1719641852
transform -1 0 1444 0 -1 2505
box -2 -3 34 103
use CLKBUF1  CLKBUF1_62
timestamp 1719641852
transform 1 0 1444 0 -1 2505
box -2 -3 74 103
use OAI22X1  OAI22X1_14
timestamp 1719641852
transform 1 0 1516 0 -1 2505
box -2 -3 42 103
use NAND2X1  NAND2X1_64
timestamp 1719641852
transform -1 0 1580 0 -1 2505
box -2 -3 26 103
use CLKBUF1  CLKBUF1_12
timestamp 1719641852
transform 1 0 1580 0 -1 2505
box -2 -3 74 103
use OAI21X1  OAI21X1_785
timestamp 1719641852
transform 1 0 1652 0 -1 2505
box -2 -3 34 103
use OAI22X1  OAI22X1_8
timestamp 1719641852
transform 1 0 1684 0 -1 2505
box -2 -3 42 103
use INVX1  INVX1_32
timestamp 1719641852
transform -1 0 1740 0 -1 2505
box -2 -3 18 103
use INVX2  INVX2_115
timestamp 1719641852
transform 1 0 1740 0 -1 2505
box -2 -3 18 103
use AOI21X1  AOI21X1_239
timestamp 1719641852
transform -1 0 1788 0 -1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_238
timestamp 1719641852
transform -1 0 1820 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_639
timestamp 1719641852
transform -1 0 1852 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_670
timestamp 1719641852
transform 1 0 1852 0 -1 2505
box -2 -3 34 103
use FILL  FILL_24_3_0
timestamp 1719641852
transform 1 0 1884 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_3_1
timestamp 1719641852
transform 1 0 1892 0 -1 2505
box -2 -3 10 103
use NAND2X1  NAND2X1_291
timestamp 1719641852
transform 1 0 1900 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_669
timestamp 1719641852
transform -1 0 1956 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_685
timestamp 1719641852
transform 1 0 1956 0 -1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_301
timestamp 1719641852
transform -1 0 2012 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_686
timestamp 1719641852
transform -1 0 2044 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_274
timestamp 1719641852
transform -1 0 2068 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_684
timestamp 1719641852
transform 1 0 2068 0 -1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_300
timestamp 1719641852
transform 1 0 2100 0 -1 2505
box -2 -3 26 103
use BUFX4  BUFX4_58
timestamp 1719641852
transform 1 0 2124 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_590
timestamp 1719641852
transform 1 0 2156 0 -1 2505
box -2 -3 34 103
use BUFX4  BUFX4_61
timestamp 1719641852
transform 1 0 2188 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_252
timestamp 1719641852
transform 1 0 2220 0 -1 2505
box -2 -3 26 103
use BUFX4  BUFX4_36
timestamp 1719641852
transform 1 0 2244 0 -1 2505
box -2 -3 34 103
use INVX1  INVX1_137
timestamp 1719641852
transform -1 0 2292 0 -1 2505
box -2 -3 18 103
use NOR2X1  NOR2X1_264
timestamp 1719641852
transform -1 0 2316 0 -1 2505
box -2 -3 26 103
use AOI21X1  AOI21X1_187
timestamp 1719641852
transform 1 0 2316 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_250
timestamp 1719641852
transform 1 0 2348 0 -1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_263
timestamp 1719641852
transform 1 0 2372 0 -1 2505
box -2 -3 26 103
use FILL  FILL_24_4_0
timestamp 1719641852
transform -1 0 2404 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_4_1
timestamp 1719641852
transform -1 0 2412 0 -1 2505
box -2 -3 10 103
use INVX1  INVX1_136
timestamp 1719641852
transform -1 0 2428 0 -1 2505
box -2 -3 18 103
use INVX2  INVX2_79
timestamp 1719641852
transform 1 0 2428 0 -1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_482
timestamp 1719641852
transform 1 0 2444 0 -1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_168
timestamp 1719641852
transform -1 0 2508 0 -1 2505
box -2 -3 34 103
use INVX2  INVX2_104
timestamp 1719641852
transform 1 0 2508 0 -1 2505
box -2 -3 18 103
use DFFSR  DFFSR_198
timestamp 1719641852
transform -1 0 2700 0 -1 2505
box -2 -3 178 103
use OAI21X1  OAI21X1_431
timestamp 1719641852
transform -1 0 2732 0 -1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_253
timestamp 1719641852
transform 1 0 2732 0 -1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_251
timestamp 1719641852
transform 1 0 2756 0 -1 2505
box -2 -3 26 103
use AOI21X1  AOI21X1_161
timestamp 1719641852
transform 1 0 2780 0 -1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_145
timestamp 1719641852
transform 1 0 2812 0 -1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_141
timestamp 1719641852
transform -1 0 2876 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_376
timestamp 1719641852
transform -1 0 2908 0 -1 2505
box -2 -3 34 103
use FILL  FILL_24_5_0
timestamp 1719641852
transform -1 0 2916 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_5_1
timestamp 1719641852
transform -1 0 2924 0 -1 2505
box -2 -3 10 103
use AOI21X1  AOI21X1_120
timestamp 1719641852
transform -1 0 2956 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_310
timestamp 1719641852
transform 1 0 2956 0 -1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_96
timestamp 1719641852
transform 1 0 2988 0 -1 2505
box -2 -3 34 103
use NAND3X1  NAND3X1_207
timestamp 1719641852
transform 1 0 3020 0 -1 2505
box -2 -3 34 103
use INVX2  INVX2_55
timestamp 1719641852
transform -1 0 3068 0 -1 2505
box -2 -3 18 103
use NAND2X1  NAND2X1_194
timestamp 1719641852
transform 1 0 3068 0 -1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_167
timestamp 1719641852
transform 1 0 3092 0 -1 2505
box -2 -3 26 103
use AOI21X1  AOI21X1_55
timestamp 1719641852
transform 1 0 3116 0 -1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_174
timestamp 1719641852
transform 1 0 3148 0 -1 2505
box -2 -3 26 103
use AOI21X1  AOI21X1_71
timestamp 1719641852
transform 1 0 3172 0 -1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_69
timestamp 1719641852
transform 1 0 3204 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_154
timestamp 1719641852
transform 1 0 3236 0 -1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_172
timestamp 1719641852
transform 1 0 3260 0 -1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_151
timestamp 1719641852
transform 1 0 3284 0 -1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_155
timestamp 1719641852
transform 1 0 3308 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_255
timestamp 1719641852
transform 1 0 3332 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_253
timestamp 1719641852
transform 1 0 3364 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_94
timestamp 1719641852
transform 1 0 3396 0 -1 2505
box -2 -3 26 103
use FILL  FILL_24_6_0
timestamp 1719641852
transform 1 0 3420 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_6_1
timestamp 1719641852
transform 1 0 3428 0 -1 2505
box -2 -3 10 103
use OAI21X1  OAI21X1_217
timestamp 1719641852
transform 1 0 3436 0 -1 2505
box -2 -3 34 103
use NAND3X1  NAND3X1_156
timestamp 1719641852
transform -1 0 3500 0 -1 2505
box -2 -3 34 103
use NAND3X1  NAND3X1_120
timestamp 1719641852
transform -1 0 3532 0 -1 2505
box -2 -3 34 103
use NAND3X1  NAND3X1_134
timestamp 1719641852
transform -1 0 3564 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_116
timestamp 1719641852
transform 1 0 3564 0 -1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_114
timestamp 1719641852
transform 1 0 3588 0 -1 2505
box -2 -3 26 103
use BUFX4  BUFX4_247
timestamp 1719641852
transform 1 0 3612 0 -1 2505
box -2 -3 34 103
use XOR2X1  XOR2X1_2
timestamp 1719641852
transform 1 0 3644 0 -1 2505
box -2 -3 58 103
use XNOR2X1  XNOR2X1_6
timestamp 1719641852
transform 1 0 3700 0 -1 2505
box -2 -3 58 103
use FILL  FILL_25_1
timestamp 1719641852
transform -1 0 3764 0 -1 2505
box -2 -3 10 103
use FILL  FILL_25_2
timestamp 1719641852
transform -1 0 3772 0 -1 2505
box -2 -3 10 103
use FILL  FILL_25_3
timestamp 1719641852
transform -1 0 3780 0 -1 2505
box -2 -3 10 103
use BUFX2  BUFX2_40
timestamp 1719641852
transform -1 0 28 0 1 2505
box -2 -3 26 103
use DFFSR  DFFSR_69
timestamp 1719641852
transform -1 0 204 0 1 2505
box -2 -3 178 103
use DFFSR  DFFSR_15
timestamp 1719641852
transform -1 0 380 0 1 2505
box -2 -3 178 103
use FILL  FILL_25_0_0
timestamp 1719641852
transform -1 0 388 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_0_1
timestamp 1719641852
transform -1 0 396 0 1 2505
box -2 -3 10 103
use DFFSR  DFFSR_52
timestamp 1719641852
transform -1 0 572 0 1 2505
box -2 -3 178 103
use OAI21X1  OAI21X1_121
timestamp 1719641852
transform -1 0 604 0 1 2505
box -2 -3 34 103
use INVX2  INVX2_36
timestamp 1719641852
transform 1 0 604 0 1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_64
timestamp 1719641852
transform 1 0 620 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_110
timestamp 1719641852
transform -1 0 684 0 1 2505
box -2 -3 34 103
use NAND3X1  NAND3X1_34
timestamp 1719641852
transform 1 0 684 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_63
timestamp 1719641852
transform -1 0 748 0 1 2505
box -2 -3 34 103
use NAND3X1  NAND3X1_30
timestamp 1719641852
transform 1 0 748 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_55
timestamp 1719641852
transform 1 0 780 0 1 2505
box -2 -3 34 103
use NAND3X1  NAND3X1_31
timestamp 1719641852
transform 1 0 812 0 1 2505
box -2 -3 34 103
use FILL  FILL_25_1_0
timestamp 1719641852
transform 1 0 844 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_1_1
timestamp 1719641852
transform 1 0 852 0 1 2505
box -2 -3 10 103
use OAI21X1  OAI21X1_57
timestamp 1719641852
transform 1 0 860 0 1 2505
box -2 -3 34 103
use BUFX4  BUFX4_200
timestamp 1719641852
transform -1 0 924 0 1 2505
box -2 -3 34 103
use BUFX4  BUFX4_79
timestamp 1719641852
transform -1 0 956 0 1 2505
box -2 -3 34 103
use BUFX4  BUFX4_80
timestamp 1719641852
transform 1 0 956 0 1 2505
box -2 -3 34 103
use BUFX4  BUFX4_86
timestamp 1719641852
transform 1 0 988 0 1 2505
box -2 -3 34 103
use INVX8  INVX8_2
timestamp 1719641852
transform -1 0 1060 0 1 2505
box -2 -3 42 103
use NAND2X1  NAND2X1_28
timestamp 1719641852
transform 1 0 1060 0 1 2505
box -2 -3 26 103
use INVX1  INVX1_26
timestamp 1719641852
transform -1 0 1100 0 1 2505
box -2 -3 18 103
use NAND2X1  NAND2X1_239
timestamp 1719641852
transform 1 0 1100 0 1 2505
box -2 -3 26 103
use OAI22X1  OAI22X1_18
timestamp 1719641852
transform 1 0 1124 0 1 2505
box -2 -3 42 103
use OAI21X1  OAI21X1_265
timestamp 1719641852
transform -1 0 1196 0 1 2505
box -2 -3 34 103
use OAI22X1  OAI22X1_15
timestamp 1719641852
transform -1 0 1236 0 1 2505
box -2 -3 42 103
use OAI22X1  OAI22X1_9
timestamp 1719641852
transform -1 0 1276 0 1 2505
box -2 -3 42 103
use NAND2X1  NAND2X1_243
timestamp 1719641852
transform -1 0 1300 0 1 2505
box -2 -3 26 103
use FILL  FILL_25_2_0
timestamp 1719641852
transform 1 0 1300 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_2_1
timestamp 1719641852
transform 1 0 1308 0 1 2505
box -2 -3 10 103
use DFFSR  DFFSR_139
timestamp 1719641852
transform 1 0 1316 0 1 2505
box -2 -3 178 103
use INVX2  INVX2_131
timestamp 1719641852
transform 1 0 1492 0 1 2505
box -2 -3 18 103
use NAND2X1  NAND2X1_67
timestamp 1719641852
transform 1 0 1508 0 1 2505
box -2 -3 26 103
use NAND3X1  NAND3X1_90
timestamp 1719641852
transform -1 0 1564 0 1 2505
box -2 -3 34 103
use DFFSR  DFFSR_151
timestamp 1719641852
transform 1 0 1564 0 1 2505
box -2 -3 178 103
use NOR2X1  NOR2X1_292
timestamp 1719641852
transform 1 0 1740 0 1 2505
box -2 -3 26 103
use AOI22X1  AOI22X1_15
timestamp 1719641852
transform 1 0 1764 0 1 2505
box -2 -3 42 103
use NAND3X1  NAND3X1_93
timestamp 1719641852
transform -1 0 1836 0 1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_202
timestamp 1719641852
transform -1 0 1868 0 1 2505
box -2 -3 34 103
use FILL  FILL_25_3_0
timestamp 1719641852
transform -1 0 1876 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_3_1
timestamp 1719641852
transform -1 0 1884 0 1 2505
box -2 -3 10 103
use OAI21X1  OAI21X1_592
timestamp 1719641852
transform -1 0 1916 0 1 2505
box -2 -3 34 103
use INVX2  INVX2_80
timestamp 1719641852
transform 1 0 1916 0 1 2505
box -2 -3 18 103
use DFFSR  DFFSR_134
timestamp 1719641852
transform -1 0 2108 0 1 2505
box -2 -3 178 103
use NAND2X1  NAND2X1_299
timestamp 1719641852
transform -1 0 2132 0 1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_309
timestamp 1719641852
transform -1 0 2156 0 1 2505
box -2 -3 26 103
use DFFSR  DFFSR_181
timestamp 1719641852
transform -1 0 2332 0 1 2505
box -2 -3 178 103
use OAI21X1  OAI21X1_549
timestamp 1719641852
transform 1 0 2332 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_552
timestamp 1719641852
transform -1 0 2396 0 1 2505
box -2 -3 34 103
use FILL  FILL_25_4_0
timestamp 1719641852
transform 1 0 2396 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_4_1
timestamp 1719641852
transform 1 0 2404 0 1 2505
box -2 -3 10 103
use OAI21X1  OAI21X1_597
timestamp 1719641852
transform 1 0 2412 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_551
timestamp 1719641852
transform -1 0 2476 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_550
timestamp 1719641852
transform -1 0 2508 0 1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_186
timestamp 1719641852
transform 1 0 2508 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_544
timestamp 1719641852
transform 1 0 2540 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_607
timestamp 1719641852
transform 1 0 2572 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_485
timestamp 1719641852
transform -1 0 2636 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_484
timestamp 1719641852
transform 1 0 2636 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_483
timestamp 1719641852
transform -1 0 2700 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_377
timestamp 1719641852
transform -1 0 2732 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_491
timestamp 1719641852
transform 1 0 2732 0 1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_170
timestamp 1719641852
transform -1 0 2796 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_465
timestamp 1719641852
transform 1 0 2796 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_378
timestamp 1719641852
transform 1 0 2828 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_428
timestamp 1719641852
transform -1 0 2892 0 1 2505
box -2 -3 34 103
use INVX2  INVX2_148
timestamp 1719641852
transform 1 0 2892 0 1 2505
box -2 -3 18 103
use FILL  FILL_25_5_0
timestamp 1719641852
transform 1 0 2908 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_5_1
timestamp 1719641852
transform 1 0 2916 0 1 2505
box -2 -3 10 103
use OAI21X1  OAI21X1_379
timestamp 1719641852
transform 1 0 2924 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_375
timestamp 1719641852
transform -1 0 2988 0 1 2505
box -2 -3 34 103
use INVX2  INVX2_73
timestamp 1719641852
transform -1 0 3004 0 1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_311
timestamp 1719641852
transform 1 0 3004 0 1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_72
timestamp 1719641852
transform 1 0 3036 0 1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_152
timestamp 1719641852
transform 1 0 3068 0 1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_154
timestamp 1719641852
transform 1 0 3092 0 1 2505
box -2 -3 26 103
use AOI22X1  AOI22X1_38
timestamp 1719641852
transform 1 0 3116 0 1 2505
box -2 -3 42 103
use INVX1  INVX1_118
timestamp 1719641852
transform 1 0 3156 0 1 2505
box -2 -3 18 103
use AOI22X1  AOI22X1_48
timestamp 1719641852
transform -1 0 3212 0 1 2505
box -2 -3 42 103
use NAND2X1  NAND2X1_173
timestamp 1719641852
transform -1 0 3236 0 1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_171
timestamp 1719641852
transform 1 0 3236 0 1 2505
box -2 -3 26 103
use AOI22X1  AOI22X1_47
timestamp 1719641852
transform 1 0 3260 0 1 2505
box -2 -3 42 103
use NAND2X1  NAND2X1_175
timestamp 1719641852
transform 1 0 3300 0 1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_150
timestamp 1719641852
transform 1 0 3324 0 1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_153
timestamp 1719641852
transform 1 0 3348 0 1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_254
timestamp 1719641852
transform 1 0 3372 0 1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_93
timestamp 1719641852
transform 1 0 3404 0 1 2505
box -2 -3 26 103
use FILL  FILL_25_6_0
timestamp 1719641852
transform -1 0 3436 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_6_1
timestamp 1719641852
transform -1 0 3444 0 1 2505
box -2 -3 10 103
use NOR2X1  NOR2X1_91
timestamp 1719641852
transform -1 0 3468 0 1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_216
timestamp 1719641852
transform 1 0 3468 0 1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_121
timestamp 1719641852
transform 1 0 3500 0 1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_122
timestamp 1719641852
transform 1 0 3524 0 1 2505
box -2 -3 26 103
use BUFX4  BUFX4_217
timestamp 1719641852
transform -1 0 3580 0 1 2505
box -2 -3 34 103
use BUFX4  BUFX4_45
timestamp 1719641852
transform -1 0 3612 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_183
timestamp 1719641852
transform -1 0 3644 0 1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_109
timestamp 1719641852
transform -1 0 3668 0 1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_202
timestamp 1719641852
transform 1 0 3668 0 1 2505
box -2 -3 34 103
use INVX1  INVX1_90
timestamp 1719641852
transform 1 0 3700 0 1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_186
timestamp 1719641852
transform 1 0 3716 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_201
timestamp 1719641852
transform 1 0 3748 0 1 2505
box -2 -3 34 103
use CLKBUF1  CLKBUF1_41
timestamp 1719641852
transform 1 0 4 0 -1 2705
box -2 -3 74 103
use CLKBUF1  CLKBUF1_35
timestamp 1719641852
transform 1 0 76 0 -1 2705
box -2 -3 74 103
use DFFSR  DFFSR_48
timestamp 1719641852
transform 1 0 148 0 -1 2705
box -2 -3 178 103
use INVX2  INVX2_12
timestamp 1719641852
transform 1 0 324 0 -1 2705
box -2 -3 18 103
use FILL  FILL_26_0_0
timestamp 1719641852
transform 1 0 340 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_0_1
timestamp 1719641852
transform 1 0 348 0 -1 2705
box -2 -3 10 103
use INVX2  INVX2_32
timestamp 1719641852
transform 1 0 356 0 -1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_56
timestamp 1719641852
transform -1 0 404 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_113
timestamp 1719641852
transform -1 0 436 0 -1 2705
box -2 -3 34 103
use INVX2  INVX2_35
timestamp 1719641852
transform 1 0 436 0 -1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_58
timestamp 1719641852
transform 1 0 452 0 -1 2705
box -2 -3 34 103
use NAND3X1  NAND3X1_60
timestamp 1719641852
transform -1 0 516 0 -1 2705
box -2 -3 34 103
use AND2X2  AND2X2_2
timestamp 1719641852
transform -1 0 548 0 -1 2705
box -2 -3 34 103
use NAND3X1  NAND3X1_64
timestamp 1719641852
transform -1 0 580 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_120
timestamp 1719641852
transform -1 0 612 0 -1 2705
box -2 -3 34 103
use OAI22X1  OAI22X1_13
timestamp 1719641852
transform -1 0 652 0 -1 2705
box -2 -3 42 103
use INVX1  INVX1_25
timestamp 1719641852
transform -1 0 668 0 -1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_92
timestamp 1719641852
transform 1 0 668 0 -1 2705
box -2 -3 34 103
use OAI22X1  OAI22X1_6
timestamp 1719641852
transform 1 0 700 0 -1 2705
box -2 -3 42 103
use NOR2X1  NOR2X1_6
timestamp 1719641852
transform -1 0 764 0 -1 2705
box -2 -3 26 103
use OAI22X1  OAI22X1_5
timestamp 1719641852
transform 1 0 764 0 -1 2705
box -2 -3 42 103
use OAI22X1  OAI22X1_3
timestamp 1719641852
transform 1 0 804 0 -1 2705
box -2 -3 42 103
use NAND2X1  NAND2X1_31
timestamp 1719641852
transform -1 0 868 0 -1 2705
box -2 -3 26 103
use FILL  FILL_26_1_0
timestamp 1719641852
transform -1 0 876 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_1_1
timestamp 1719641852
transform -1 0 884 0 -1 2705
box -2 -3 10 103
use NAND3X1  NAND3X1_77
timestamp 1719641852
transform -1 0 916 0 -1 2705
box -2 -3 34 103
use OAI22X1  OAI22X1_2
timestamp 1719641852
transform 1 0 916 0 -1 2705
box -2 -3 42 103
use NOR2X1  NOR2X1_2
timestamp 1719641852
transform -1 0 980 0 -1 2705
box -2 -3 26 103
use OAI22X1  OAI22X1_1
timestamp 1719641852
transform 1 0 980 0 -1 2705
box -2 -3 42 103
use INVX1  INVX1_30
timestamp 1719641852
transform -1 0 1036 0 -1 2705
box -2 -3 18 103
use INVX1  INVX1_31
timestamp 1719641852
transform -1 0 1052 0 -1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_84
timestamp 1719641852
transform -1 0 1084 0 -1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_9
timestamp 1719641852
transform 1 0 1084 0 -1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_44
timestamp 1719641852
transform -1 0 1132 0 -1 2705
box -2 -3 26 103
use DFFSR  DFFSR_244
timestamp 1719641852
transform -1 0 1308 0 -1 2705
box -2 -3 178 103
use FILL  FILL_26_2_0
timestamp 1719641852
transform 1 0 1308 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_2_1
timestamp 1719641852
transform 1 0 1316 0 -1 2705
box -2 -3 10 103
use DFFSR  DFFSR_169
timestamp 1719641852
transform 1 0 1324 0 -1 2705
box -2 -3 178 103
use INVX2  INVX2_163
timestamp 1719641852
transform 1 0 1500 0 -1 2705
box -2 -3 18 103
use INVX1  INVX1_38
timestamp 1719641852
transform -1 0 1532 0 -1 2705
box -2 -3 18 103
use NOR2X1  NOR2X1_275
timestamp 1719641852
transform 1 0 1532 0 -1 2705
box -2 -3 26 103
use AOI21X1  AOI21X1_203
timestamp 1719641852
transform -1 0 1588 0 -1 2705
box -2 -3 34 103
use INVX2  INVX2_76
timestamp 1719641852
transform 1 0 1588 0 -1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_641
timestamp 1719641852
transform 1 0 1604 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_642
timestamp 1719641852
transform -1 0 1668 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_591
timestamp 1719641852
transform -1 0 1700 0 -1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_201
timestamp 1719641852
transform 1 0 1700 0 -1 2705
box -2 -3 34 103
use OR2X2  OR2X2_16
timestamp 1719641852
transform -1 0 1764 0 -1 2705
box -2 -3 34 103
use INVX2  INVX2_56
timestamp 1719641852
transform -1 0 1780 0 -1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_640
timestamp 1719641852
transform -1 0 1812 0 -1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_323
timestamp 1719641852
transform 1 0 1812 0 -1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_322
timestamp 1719641852
transform 1 0 1836 0 -1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_726
timestamp 1719641852
transform -1 0 1892 0 -1 2705
box -2 -3 34 103
use FILL  FILL_26_3_0
timestamp 1719641852
transform -1 0 1900 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_3_1
timestamp 1719641852
transform -1 0 1908 0 -1 2705
box -2 -3 10 103
use DFFSR  DFFSR_182
timestamp 1719641852
transform -1 0 2084 0 -1 2705
box -2 -3 178 103
use INVX1  INVX1_27
timestamp 1719641852
transform -1 0 2100 0 -1 2705
box -2 -3 18 103
use NOR2X1  NOR2X1_293
timestamp 1719641852
transform 1 0 2100 0 -1 2705
box -2 -3 26 103
use INVX2  INVX2_159
timestamp 1719641852
transform 1 0 2124 0 -1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_548
timestamp 1719641852
transform 1 0 2140 0 -1 2705
box -2 -3 34 103
use INVX2  INVX2_146
timestamp 1719641852
transform 1 0 2172 0 -1 2705
box -2 -3 18 103
use AOI21X1  AOI21X1_169
timestamp 1719641852
transform 1 0 2188 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_487
timestamp 1719641852
transform 1 0 2220 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_543
timestamp 1719641852
transform 1 0 2252 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_547
timestamp 1719641852
transform -1 0 2316 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_546
timestamp 1719641852
transform -1 0 2348 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_545
timestamp 1719641852
transform -1 0 2380 0 -1 2705
box -2 -3 34 103
use FILL  FILL_26_4_0
timestamp 1719641852
transform 1 0 2380 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_4_1
timestamp 1719641852
transform 1 0 2388 0 -1 2705
box -2 -3 10 103
use OAI21X1  OAI21X1_481
timestamp 1719641852
transform 1 0 2396 0 -1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_280
timestamp 1719641852
transform -1 0 2452 0 -1 2705
box -2 -3 26 103
use DFFSR  DFFSR_232
timestamp 1719641852
transform -1 0 2628 0 -1 2705
box -2 -3 178 103
use INVX2  INVX2_89
timestamp 1719641852
transform 1 0 2628 0 -1 2705
box -2 -3 18 103
use NOR2X1  NOR2X1_213
timestamp 1719641852
transform 1 0 2644 0 -1 2705
box -2 -3 26 103
use AOI21X1  AOI21X1_115
timestamp 1719641852
transform -1 0 2700 0 -1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_217
timestamp 1719641852
transform 1 0 2700 0 -1 2705
box -2 -3 26 103
use AOI21X1  AOI21X1_123
timestamp 1719641852
transform -1 0 2756 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_466
timestamp 1719641852
transform -1 0 2788 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_467
timestamp 1719641852
transform 1 0 2788 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_429
timestamp 1719641852
transform -1 0 2852 0 -1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_162
timestamp 1719641852
transform 1 0 2852 0 -1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_244
timestamp 1719641852
transform -1 0 2908 0 -1 2705
box -2 -3 26 103
use FILL  FILL_26_5_0
timestamp 1719641852
transform 1 0 2908 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_5_1
timestamp 1719641852
transform 1 0 2916 0 -1 2705
box -2 -3 10 103
use NOR2X1  NOR2X1_229
timestamp 1719641852
transform 1 0 2924 0 -1 2705
box -2 -3 26 103
use INVX2  INVX2_75
timestamp 1719641852
transform 1 0 2948 0 -1 2705
box -2 -3 18 103
use DFFSR  DFFSR_202
timestamp 1719641852
transform 1 0 2964 0 -1 2705
box -2 -3 178 103
use OAI21X1  OAI21X1_295
timestamp 1719641852
transform -1 0 3172 0 -1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_97
timestamp 1719641852
transform -1 0 3204 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_293
timestamp 1719641852
transform -1 0 3236 0 -1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_152
timestamp 1719641852
transform 1 0 3236 0 -1 2705
box -2 -3 26 103
use AOI21X1  AOI21X1_70
timestamp 1719641852
transform 1 0 3260 0 -1 2705
box -2 -3 34 103
use BUFX4  BUFX4_172
timestamp 1719641852
transform -1 0 3324 0 -1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_156
timestamp 1719641852
transform 1 0 3324 0 -1 2705
box -2 -3 26 103
use NOR2X1  NOR2X1_157
timestamp 1719641852
transform 1 0 3348 0 -1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_256
timestamp 1719641852
transform 1 0 3372 0 -1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_92
timestamp 1719641852
transform 1 0 3404 0 -1 2705
box -2 -3 26 103
use FILL  FILL_26_6_0
timestamp 1719641852
transform -1 0 3436 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_6_1
timestamp 1719641852
transform -1 0 3444 0 -1 2705
box -2 -3 10 103
use NOR2X1  NOR2X1_117
timestamp 1719641852
transform -1 0 3468 0 -1 2705
box -2 -3 26 103
use NOR2X1  NOR2X1_118
timestamp 1719641852
transform -1 0 3492 0 -1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_235
timestamp 1719641852
transform 1 0 3492 0 -1 2705
box -2 -3 34 103
use NAND3X1  NAND3X1_194
timestamp 1719641852
transform -1 0 3556 0 -1 2705
box -2 -3 34 103
use NAND3X1  NAND3X1_196
timestamp 1719641852
transform 1 0 3556 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_291
timestamp 1719641852
transform -1 0 3620 0 -1 2705
box -2 -3 34 103
use INVX1  INVX1_106
timestamp 1719641852
transform -1 0 3636 0 -1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_294
timestamp 1719641852
transform 1 0 3636 0 -1 2705
box -2 -3 34 103
use INVX1  INVX1_81
timestamp 1719641852
transform 1 0 3668 0 -1 2705
box -2 -3 18 103
use NOR2X1  NOR2X1_54
timestamp 1719641852
transform -1 0 3708 0 -1 2705
box -2 -3 26 103
use INVX1  INVX1_83
timestamp 1719641852
transform 1 0 3708 0 -1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_185
timestamp 1719641852
transform 1 0 3724 0 -1 2705
box -2 -3 34 103
use FILL  FILL_27_1
timestamp 1719641852
transform -1 0 3764 0 -1 2705
box -2 -3 10 103
use FILL  FILL_27_2
timestamp 1719641852
transform -1 0 3772 0 -1 2705
box -2 -3 10 103
use FILL  FILL_27_3
timestamp 1719641852
transform -1 0 3780 0 -1 2705
box -2 -3 10 103
use BUFX2  BUFX2_58
timestamp 1719641852
transform -1 0 28 0 1 2705
box -2 -3 26 103
use DFFSR  DFFSR_87
timestamp 1719641852
transform -1 0 204 0 1 2705
box -2 -3 178 103
use DFFSR  DFFSR_4
timestamp 1719641852
transform -1 0 380 0 1 2705
box -2 -3 178 103
use FILL  FILL_27_0_0
timestamp 1719641852
transform 1 0 380 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_0_1
timestamp 1719641852
transform 1 0 388 0 1 2705
box -2 -3 10 103
use DFFSR  DFFSR_49
timestamp 1719641852
transform 1 0 396 0 1 2705
box -2 -3 178 103
use INVX2  INVX2_13
timestamp 1719641852
transform 1 0 572 0 1 2705
box -2 -3 18 103
use NAND3X1  NAND3X1_41
timestamp 1719641852
transform -1 0 620 0 1 2705
box -2 -3 34 103
use INVX2  INVX2_33
timestamp 1719641852
transform 1 0 620 0 1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_115
timestamp 1719641852
transform 1 0 636 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_93
timestamp 1719641852
transform 1 0 668 0 1 2705
box -2 -3 34 103
use NAND3X1  NAND3X1_49
timestamp 1719641852
transform 1 0 700 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_119
timestamp 1719641852
transform 1 0 732 0 1 2705
box -2 -3 34 103
use NAND3X1  NAND3X1_61
timestamp 1719641852
transform 1 0 764 0 1 2705
box -2 -3 34 103
use NAND3X1  NAND3X1_63
timestamp 1719641852
transform 1 0 796 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_114
timestamp 1719641852
transform 1 0 828 0 1 2705
box -2 -3 34 103
use FILL  FILL_27_1_0
timestamp 1719641852
transform -1 0 868 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_1_1
timestamp 1719641852
transform -1 0 876 0 1 2705
box -2 -3 10 103
use OAI21X1  OAI21X1_112
timestamp 1719641852
transform -1 0 908 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_118
timestamp 1719641852
transform -1 0 940 0 1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_29
timestamp 1719641852
transform -1 0 964 0 1 2705
box -2 -3 26 103
use NOR2X1  NOR2X1_5
timestamp 1719641852
transform 1 0 964 0 1 2705
box -2 -3 26 103
use OAI22X1  OAI22X1_4
timestamp 1719641852
transform 1 0 988 0 1 2705
box -2 -3 42 103
use BUFX4  BUFX4_85
timestamp 1719641852
transform 1 0 1028 0 1 2705
box -2 -3 34 103
use BUFX4  BUFX4_83
timestamp 1719641852
transform 1 0 1060 0 1 2705
box -2 -3 34 103
use BUFX4  BUFX4_84
timestamp 1719641852
transform 1 0 1092 0 1 2705
box -2 -3 34 103
use DFFSR  DFFSR_68
timestamp 1719641852
transform -1 0 1300 0 1 2705
box -2 -3 178 103
use AOI21X1  AOI21X1_6
timestamp 1719641852
transform -1 0 1332 0 1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_242
timestamp 1719641852
transform -1 0 1356 0 1 2705
box -2 -3 26 103
use FILL  FILL_27_2_0
timestamp 1719641852
transform 1 0 1356 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_2_1
timestamp 1719641852
transform 1 0 1364 0 1 2705
box -2 -3 10 103
use BUFX4  BUFX4_25
timestamp 1719641852
transform 1 0 1372 0 1 2705
box -2 -3 34 103
use NAND3X1  NAND3X1_71
timestamp 1719641852
transform 1 0 1404 0 1 2705
box -2 -3 34 103
use BUFX4  BUFX4_193
timestamp 1719641852
transform 1 0 1436 0 1 2705
box -2 -3 34 103
use AOI22X1  AOI22X1_10
timestamp 1719641852
transform 1 0 1468 0 1 2705
box -2 -3 42 103
use DFFSR  DFFSR_118
timestamp 1719641852
transform -1 0 1684 0 1 2705
box -2 -3 178 103
use AOI22X1  AOI22X1_14
timestamp 1719641852
transform 1 0 1684 0 1 2705
box -2 -3 42 103
use NAND3X1  NAND3X1_92
timestamp 1719641852
transform -1 0 1756 0 1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_66
timestamp 1719641852
transform -1 0 1780 0 1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_244
timestamp 1719641852
transform -1 0 1804 0 1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_280
timestamp 1719641852
transform 1 0 1804 0 1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_643
timestamp 1719641852
transform -1 0 1860 0 1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_240
timestamp 1719641852
transform -1 0 1892 0 1 2705
box -2 -3 34 103
use FILL  FILL_27_3_0
timestamp 1719641852
transform -1 0 1900 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_3_1
timestamp 1719641852
transform -1 0 1908 0 1 2705
box -2 -3 10 103
use OAI21X1  OAI21X1_728
timestamp 1719641852
transform -1 0 1940 0 1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_322
timestamp 1719641852
transform -1 0 1964 0 1 2705
box -2 -3 26 103
use INVX1  INVX1_159
timestamp 1719641852
transform 1 0 1964 0 1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_727
timestamp 1719641852
transform 1 0 1980 0 1 2705
box -2 -3 34 103
use INVX2  INVX2_74
timestamp 1719641852
transform 1 0 2012 0 1 2705
box -2 -3 18 103
use AOI22X1  AOI22X1_13
timestamp 1719641852
transform 1 0 2028 0 1 2705
box -2 -3 42 103
use DFFSR  DFFSR_197
timestamp 1719641852
transform -1 0 2244 0 1 2705
box -2 -3 178 103
use INVX2  INVX2_149
timestamp 1719641852
transform -1 0 2260 0 1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_490
timestamp 1719641852
transform -1 0 2292 0 1 2705
box -2 -3 34 103
use INVX2  INVX2_105
timestamp 1719641852
transform 1 0 2292 0 1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_489
timestamp 1719641852
transform -1 0 2340 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_488
timestamp 1719641852
transform -1 0 2372 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_554
timestamp 1719641852
transform -1 0 2404 0 1 2705
box -2 -3 34 103
use FILL  FILL_27_4_0
timestamp 1719641852
transform -1 0 2412 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_4_1
timestamp 1719641852
transform -1 0 2420 0 1 2705
box -2 -3 10 103
use AOI21X1  AOI21X1_188
timestamp 1719641852
transform -1 0 2452 0 1 2705
box -2 -3 34 103
use DFFSR  DFFSR_228
timestamp 1719641852
transform -1 0 2628 0 1 2705
box -2 -3 178 103
use OAI21X1  OAI21X1_367
timestamp 1719641852
transform -1 0 2660 0 1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_114
timestamp 1719641852
transform 1 0 2660 0 1 2705
box -2 -3 34 103
use INVX2  INVX2_102
timestamp 1719641852
transform 1 0 2692 0 1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_381
timestamp 1719641852
transform 1 0 2708 0 1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_122
timestamp 1719641852
transform 1 0 2740 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_492
timestamp 1719641852
transform -1 0 2804 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_493
timestamp 1719641852
transform 1 0 2804 0 1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_142
timestamp 1719641852
transform -1 0 2868 0 1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_143
timestamp 1719641852
transform 1 0 2868 0 1 2705
box -2 -3 34 103
use FILL  FILL_27_5_0
timestamp 1719641852
transform -1 0 2908 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_5_1
timestamp 1719641852
transform -1 0 2916 0 1 2705
box -2 -3 10 103
use DFFSR  DFFSR_214
timestamp 1719641852
transform -1 0 3092 0 1 2705
box -2 -3 178 103
use DFFSR  DFFSR_246
timestamp 1719641852
transform 1 0 3092 0 1 2705
box -2 -3 178 103
use OAI21X1  OAI21X1_284
timestamp 1719641852
transform 1 0 3268 0 1 2705
box -2 -3 34 103
use XOR2X1  XOR2X1_4
timestamp 1719641852
transform 1 0 3300 0 1 2705
box -2 -3 58 103
use NOR2X1  NOR2X1_184
timestamp 1719641852
transform -1 0 3380 0 1 2705
box -2 -3 26 103
use AOI21X1  AOI21X1_49
timestamp 1719641852
transform 1 0 3380 0 1 2705
box -2 -3 34 103
use FILL  FILL_27_6_0
timestamp 1719641852
transform 1 0 3412 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_6_1
timestamp 1719641852
transform 1 0 3420 0 1 2705
box -2 -3 10 103
use INVX2  INVX2_44
timestamp 1719641852
transform 1 0 3428 0 1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_286
timestamp 1719641852
transform 1 0 3444 0 1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_50
timestamp 1719641852
transform -1 0 3508 0 1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_42
timestamp 1719641852
transform 1 0 3508 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_184
timestamp 1719641852
transform -1 0 3572 0 1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_52
timestamp 1719641852
transform -1 0 3596 0 1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_182
timestamp 1719641852
transform -1 0 3628 0 1 2705
box -2 -3 34 103
use BUFX4  BUFX4_245
timestamp 1719641852
transform 1 0 3628 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_203
timestamp 1719641852
transform 1 0 3660 0 1 2705
box -2 -3 34 103
use NAND3X1  NAND3X1_108
timestamp 1719641852
transform 1 0 3692 0 1 2705
box -2 -3 34 103
use OR2X2  OR2X2_9
timestamp 1719641852
transform -1 0 3756 0 1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_112
timestamp 1719641852
transform -1 0 3780 0 1 2705
box -2 -3 26 103
use BUFX2  BUFX2_17
timestamp 1719641852
transform -1 0 28 0 -1 2905
box -2 -3 26 103
use BUFX2  BUFX2_6
timestamp 1719641852
transform -1 0 52 0 -1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_130
timestamp 1719641852
transform 1 0 52 0 -1 2905
box -2 -3 34 103
use BUFX4  BUFX4_95
timestamp 1719641852
transform -1 0 116 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_141
timestamp 1719641852
transform 1 0 116 0 -1 2905
box -2 -3 34 103
use CLKBUF1  CLKBUF1_64
timestamp 1719641852
transform -1 0 220 0 -1 2905
box -2 -3 74 103
use OAI21X1  OAI21X1_149
timestamp 1719641852
transform 1 0 220 0 -1 2905
box -2 -3 34 103
use DFFSR  DFFSR_51
timestamp 1719641852
transform 1 0 252 0 -1 2905
box -2 -3 178 103
use FILL  FILL_28_0_0
timestamp 1719641852
transform 1 0 428 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_0_1
timestamp 1719641852
transform 1 0 436 0 -1 2905
box -2 -3 10 103
use DFFSR  DFFSR_34
timestamp 1719641852
transform 1 0 444 0 -1 2905
box -2 -3 178 103
use INVX1  INVX1_22
timestamp 1719641852
transform 1 0 620 0 -1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_78
timestamp 1719641852
transform 1 0 636 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_81
timestamp 1719641852
transform 1 0 668 0 -1 2905
box -2 -3 34 103
use NAND3X1  NAND3X1_43
timestamp 1719641852
transform -1 0 732 0 -1 2905
box -2 -3 34 103
use INVX1  INVX1_23
timestamp 1719641852
transform -1 0 748 0 -1 2905
box -2 -3 18 103
use NAND2X1  NAND2X1_41
timestamp 1719641852
transform -1 0 772 0 -1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_80
timestamp 1719641852
transform 1 0 772 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_49
timestamp 1719641852
transform -1 0 836 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_61
timestamp 1719641852
transform -1 0 868 0 -1 2905
box -2 -3 34 103
use FILL  FILL_28_1_0
timestamp 1719641852
transform -1 0 876 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_1_1
timestamp 1719641852
transform -1 0 884 0 -1 2905
box -2 -3 10 103
use OAI21X1  OAI21X1_86
timestamp 1719641852
transform -1 0 916 0 -1 2905
box -2 -3 34 103
use BUFX4  BUFX4_16
timestamp 1719641852
transform 1 0 916 0 -1 2905
box -2 -3 34 103
use BUFX4  BUFX4_82
timestamp 1719641852
transform -1 0 980 0 -1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_39
timestamp 1719641852
transform -1 0 1004 0 -1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_90
timestamp 1719641852
transform -1 0 1036 0 -1 2905
box -2 -3 34 103
use NAND3X1  NAND3X1_45
timestamp 1719641852
transform -1 0 1068 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_85
timestamp 1719641852
transform -1 0 1100 0 -1 2905
box -2 -3 34 103
use DFFSR  DFFSR_36
timestamp 1719641852
transform 1 0 1100 0 -1 2905
box -2 -3 178 103
use INVX2  INVX2_19
timestamp 1719641852
transform -1 0 1292 0 -1 2905
box -2 -3 18 103
use NAND2X1  NAND2X1_25
timestamp 1719641852
transform -1 0 1316 0 -1 2905
box -2 -3 26 103
use NAND3X1  NAND3X1_72
timestamp 1719641852
transform -1 0 1348 0 -1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_3
timestamp 1719641852
transform -1 0 1380 0 -1 2905
box -2 -3 34 103
use FILL  FILL_28_2_0
timestamp 1719641852
transform -1 0 1388 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_2_1
timestamp 1719641852
transform -1 0 1396 0 -1 2905
box -2 -3 10 103
use NAND2X1  NAND2X1_38
timestamp 1719641852
transform -1 0 1420 0 -1 2905
box -2 -3 26 103
use AOI21X1  AOI21X1_2
timestamp 1719641852
transform -1 0 1452 0 -1 2905
box -2 -3 34 103
use NAND3X1  NAND3X1_73
timestamp 1719641852
transform 1 0 1452 0 -1 2905
box -2 -3 34 103
use INVX1  INVX1_29
timestamp 1719641852
transform -1 0 1500 0 -1 2905
box -2 -3 18 103
use INVX2  INVX2_18
timestamp 1719641852
transform -1 0 1516 0 -1 2905
box -2 -3 18 103
use DFFSR  DFFSR_150
timestamp 1719641852
transform -1 0 1692 0 -1 2905
box -2 -3 178 103
use AOI22X1  AOI22X1_5
timestamp 1719641852
transform 1 0 1692 0 -1 2905
box -2 -3 42 103
use BUFX4  BUFX4_246
timestamp 1719641852
transform -1 0 1764 0 -1 2905
box -2 -3 34 103
use DFFSR  DFFSR_138
timestamp 1719641852
transform -1 0 1940 0 -1 2905
box -2 -3 178 103
use FILL  FILL_28_3_0
timestamp 1719641852
transform -1 0 1948 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_3_1
timestamp 1719641852
transform -1 0 1956 0 -1 2905
box -2 -3 10 103
use BUFX4  BUFX4_204
timestamp 1719641852
transform -1 0 1988 0 -1 2905
box -2 -3 34 103
use BUFX4  BUFX4_211
timestamp 1719641852
transform 1 0 1988 0 -1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_277
timestamp 1719641852
transform 1 0 2020 0 -1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_635
timestamp 1719641852
transform -1 0 2076 0 -1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_290
timestamp 1719641852
transform -1 0 2100 0 -1 2905
box -2 -3 26 103
use AOI21X1  AOI21X1_233
timestamp 1719641852
transform 1 0 2100 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_632
timestamp 1719641852
transform 1 0 2132 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_634
timestamp 1719641852
transform -1 0 2196 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_633
timestamp 1719641852
transform -1 0 2228 0 -1 2905
box -2 -3 34 103
use BUFX4  BUFX4_121
timestamp 1719641852
transform -1 0 2260 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_486
timestamp 1719641852
transform -1 0 2292 0 -1 2905
box -2 -3 34 103
use INVX2  INVX2_106
timestamp 1719641852
transform 1 0 2292 0 -1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_602
timestamp 1719641852
transform -1 0 2340 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_556
timestamp 1719641852
transform -1 0 2372 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_555
timestamp 1719641852
transform -1 0 2404 0 -1 2905
box -2 -3 34 103
use FILL  FILL_28_4_0
timestamp 1719641852
transform 1 0 2404 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_4_1
timestamp 1719641852
transform 1 0 2412 0 -1 2905
box -2 -3 10 103
use NOR2X1  NOR2X1_295
timestamp 1719641852
transform 1 0 2420 0 -1 2905
box -2 -3 26 103
use BUFX4  BUFX4_122
timestamp 1719641852
transform 1 0 2444 0 -1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_302
timestamp 1719641852
transform 1 0 2476 0 -1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_687
timestamp 1719641852
transform -1 0 2532 0 -1 2905
box -2 -3 34 103
use INVX1  INVX1_100
timestamp 1719641852
transform -1 0 2548 0 -1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_599
timestamp 1719641852
transform -1 0 2580 0 -1 2905
box -2 -3 34 103
use INVX2  INVX2_78
timestamp 1719641852
transform 1 0 2580 0 -1 2905
box -2 -3 18 103
use AOI21X1  AOI21X1_210
timestamp 1719641852
transform 1 0 2596 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_598
timestamp 1719641852
transform 1 0 2628 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_715
timestamp 1719641852
transform -1 0 2692 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_729
timestamp 1719641852
transform -1 0 2724 0 -1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_254
timestamp 1719641852
transform -1 0 2748 0 -1 2905
box -2 -3 26 103
use AOI21X1  AOI21X1_171
timestamp 1719641852
transform -1 0 2780 0 -1 2905
box -2 -3 34 103
use INVX2  INVX2_101
timestamp 1719641852
transform 1 0 2780 0 -1 2905
box -2 -3 18 103
use INVX1  INVX1_102
timestamp 1719641852
transform -1 0 2812 0 -1 2905
box -2 -3 18 103
use DFFSR  DFFSR_229
timestamp 1719641852
transform -1 0 2988 0 -1 2905
box -2 -3 178 103
use FILL  FILL_28_5_0
timestamp 1719641852
transform 1 0 2988 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_5_1
timestamp 1719641852
transform 1 0 2996 0 -1 2905
box -2 -3 10 103
use INVX1  INVX1_99
timestamp 1719641852
transform 1 0 3004 0 -1 2905
box -2 -3 18 103
use NAND3X1  NAND3X1_200
timestamp 1719641852
transform 1 0 3020 0 -1 2905
box -2 -3 34 103
use NAND3X1  NAND3X1_201
timestamp 1719641852
transform 1 0 3052 0 -1 2905
box -2 -3 34 103
use NAND3X1  NAND3X1_199
timestamp 1719641852
transform 1 0 3084 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_791
timestamp 1719641852
transform 1 0 3116 0 -1 2905
box -2 -3 34 103
use XNOR2X1  XNOR2X1_12
timestamp 1719641852
transform -1 0 3204 0 -1 2905
box -2 -3 58 103
use XNOR2X1  XNOR2X1_7
timestamp 1719641852
transform -1 0 3260 0 -1 2905
box -2 -3 58 103
use AOI21X1  AOI21X1_34
timestamp 1719641852
transform -1 0 3292 0 -1 2905
box -2 -3 34 103
use OR2X2  OR2X2_10
timestamp 1719641852
transform -1 0 3324 0 -1 2905
box -2 -3 34 103
use NAND3X1  NAND3X1_195
timestamp 1719641852
transform 1 0 3324 0 -1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_181
timestamp 1719641852
transform -1 0 3380 0 -1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_285
timestamp 1719641852
transform 1 0 3380 0 -1 2905
box -2 -3 34 103
use FILL  FILL_28_6_0
timestamp 1719641852
transform 1 0 3412 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_6_1
timestamp 1719641852
transform 1 0 3420 0 -1 2905
box -2 -3 10 103
use INVX1  INVX1_104
timestamp 1719641852
transform 1 0 3428 0 -1 2905
box -2 -3 18 103
use NAND2X1  NAND2X1_131
timestamp 1719641852
transform 1 0 3444 0 -1 2905
box -2 -3 26 103
use XNOR2X1  XNOR2X1_3
timestamp 1719641852
transform -1 0 3524 0 -1 2905
box -2 -3 58 103
use NAND2X1  NAND2X1_149
timestamp 1719641852
transform 1 0 3524 0 -1 2905
box -2 -3 26 103
use BUFX4  BUFX4_248
timestamp 1719641852
transform 1 0 3548 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_287
timestamp 1719641852
transform 1 0 3580 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_289
timestamp 1719641852
transform -1 0 3644 0 -1 2905
box -2 -3 34 103
use INVX1  INVX1_115
timestamp 1719641852
transform -1 0 3660 0 -1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_197
timestamp 1719641852
transform 1 0 3660 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_196
timestamp 1719641852
transform -1 0 3724 0 -1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_63
timestamp 1719641852
transform 1 0 3724 0 -1 2905
box -2 -3 26 103
use NOR2X1  NOR2X1_64
timestamp 1719641852
transform -1 0 3772 0 -1 2905
box -2 -3 26 103
use FILL  FILL_29_1
timestamp 1719641852
transform -1 0 3780 0 -1 2905
box -2 -3 10 103
use BUFX2  BUFX2_25
timestamp 1719641852
transform -1 0 28 0 1 2905
box -2 -3 26 103
use CLKBUF1  CLKBUF1_7
timestamp 1719641852
transform 1 0 28 0 1 2905
box -2 -3 74 103
use CLKBUF1  CLKBUF1_9
timestamp 1719641852
transform 1 0 100 0 1 2905
box -2 -3 74 103
use CLKBUF1  CLKBUF1_18
timestamp 1719641852
transform 1 0 172 0 1 2905
box -2 -3 74 103
use CLKBUF1  CLKBUF1_3
timestamp 1719641852
transform 1 0 244 0 1 2905
box -2 -3 74 103
use FILL  FILL_29_0_0
timestamp 1719641852
transform 1 0 316 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_0_1
timestamp 1719641852
transform 1 0 324 0 1 2905
box -2 -3 10 103
use DFFSR  DFFSR_5
timestamp 1719641852
transform 1 0 332 0 1 2905
box -2 -3 178 103
use OAI21X1  OAI21X1_79
timestamp 1719641852
transform -1 0 540 0 1 2905
box -2 -3 34 103
use NAND3X1  NAND3X1_42
timestamp 1719641852
transform -1 0 572 0 1 2905
box -2 -3 34 103
use BUFX4  BUFX4_15
timestamp 1719641852
transform -1 0 604 0 1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_53
timestamp 1719641852
transform 1 0 604 0 1 2905
box -2 -3 34 103
use NAND3X1  NAND3X1_29
timestamp 1719641852
transform 1 0 636 0 1 2905
box -2 -3 34 103
use NAND3X1  NAND3X1_33
timestamp 1719641852
transform -1 0 700 0 1 2905
box -2 -3 34 103
use BUFX4  BUFX4_24
timestamp 1719641852
transform -1 0 732 0 1 2905
box -2 -3 34 103
use NAND3X1  NAND3X1_46
timestamp 1719641852
transform -1 0 764 0 1 2905
box -2 -3 34 103
use BUFX4  BUFX4_19
timestamp 1719641852
transform 1 0 764 0 1 2905
box -2 -3 34 103
use NAND3X1  NAND3X1_44
timestamp 1719641852
transform -1 0 828 0 1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_82
timestamp 1719641852
transform -1 0 860 0 1 2905
box -2 -3 34 103
use FILL  FILL_29_1_0
timestamp 1719641852
transform 1 0 860 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_1_1
timestamp 1719641852
transform 1 0 868 0 1 2905
box -2 -3 10 103
use NAND2X1  NAND2X1_27
timestamp 1719641852
transform 1 0 876 0 1 2905
box -2 -3 26 103
use NAND3X1  NAND3X1_47
timestamp 1719641852
transform -1 0 932 0 1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_88
timestamp 1719641852
transform -1 0 964 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_30
timestamp 1719641852
transform -1 0 988 0 1 2905
box -2 -3 26 103
use NAND3X1  NAND3X1_48
timestamp 1719641852
transform -1 0 1020 0 1 2905
box -2 -3 34 103
use DFFSR  DFFSR_19
timestamp 1719641852
transform 1 0 1020 0 1 2905
box -2 -3 178 103
use OAI21X1  OAI21X1_22
timestamp 1719641852
transform 1 0 1196 0 1 2905
box -2 -3 34 103
use INVX1  INVX1_11
timestamp 1719641852
transform 1 0 1228 0 1 2905
box -2 -3 18 103
use BUFX4  BUFX4_26
timestamp 1719641852
transform 1 0 1244 0 1 2905
box -2 -3 34 103
use NAND3X1  NAND3X1_13
timestamp 1719641852
transform 1 0 1276 0 1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_21
timestamp 1719641852
transform 1 0 1308 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_11
timestamp 1719641852
transform 1 0 1340 0 1 2905
box -2 -3 26 103
use FILL  FILL_29_2_0
timestamp 1719641852
transform -1 0 1372 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_2_1
timestamp 1719641852
transform -1 0 1380 0 1 2905
box -2 -3 10 103
use NAND2X1  NAND2X1_40
timestamp 1719641852
transform -1 0 1404 0 1 2905
box -2 -3 26 103
use BUFX4  BUFX4_126
timestamp 1719641852
transform 1 0 1404 0 1 2905
box -2 -3 34 103
use AOI22X1  AOI22X1_12
timestamp 1719641852
transform -1 0 1476 0 1 2905
box -2 -3 42 103
use NAND3X1  NAND3X1_69
timestamp 1719641852
transform 1 0 1476 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_222
timestamp 1719641852
transform 1 0 1508 0 1 2905
box -2 -3 26 103
use AOI22X1  AOI22X1_4
timestamp 1719641852
transform 1 0 1532 0 1 2905
box -2 -3 42 103
use NAND3X1  NAND3X1_87
timestamp 1719641852
transform -1 0 1604 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_61
timestamp 1719641852
transform -1 0 1628 0 1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_330
timestamp 1719641852
transform -1 0 1652 0 1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_224
timestamp 1719641852
transform 1 0 1652 0 1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_62
timestamp 1719641852
transform -1 0 1700 0 1 2905
box -2 -3 26 103
use NAND3X1  NAND3X1_88
timestamp 1719641852
transform -1 0 1732 0 1 2905
box -2 -3 34 103
use DFFSR  DFFSR_153
timestamp 1719641852
transform -1 0 1908 0 1 2905
box -2 -3 178 103
use FILL  FILL_29_3_0
timestamp 1719641852
transform 1 0 1908 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_3_1
timestamp 1719641852
transform 1 0 1916 0 1 2905
box -2 -3 10 103
use BUFX4  BUFX4_114
timestamp 1719641852
transform 1 0 1924 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_240
timestamp 1719641852
transform 1 0 1956 0 1 2905
box -2 -3 26 103
use AOI22X1  AOI22X1_3
timestamp 1719641852
transform -1 0 2020 0 1 2905
box -2 -3 42 103
use OAI21X1  OAI21X1_553
timestamp 1719641852
transform 1 0 2020 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_247
timestamp 1719641852
transform -1 0 2076 0 1 2905
box -2 -3 26 103
use BUFX4  BUFX4_113
timestamp 1719641852
transform 1 0 2076 0 1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_557
timestamp 1719641852
transform -1 0 2140 0 1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_688
timestamp 1719641852
transform -1 0 2172 0 1 2905
box -2 -3 34 103
use INVX1  INVX1_152
timestamp 1719641852
transform -1 0 2188 0 1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_689
timestamp 1719641852
transform 1 0 2188 0 1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_311
timestamp 1719641852
transform 1 0 2220 0 1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_303
timestamp 1719641852
transform 1 0 2244 0 1 2905
box -2 -3 26 103
use AOI22X1  AOI22X1_6
timestamp 1719641852
transform -1 0 2308 0 1 2905
box -2 -3 42 103
use AOI22X1  AOI22X1_1
timestamp 1719641852
transform 1 0 2308 0 1 2905
box -2 -3 42 103
use NOR2X1  NOR2X1_294
timestamp 1719641852
transform -1 0 2372 0 1 2905
box -2 -3 26 103
use AOI21X1  AOI21X1_241
timestamp 1719641852
transform 1 0 2372 0 1 2905
box -2 -3 34 103
use FILL  FILL_29_4_0
timestamp 1719641852
transform 1 0 2404 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_4_1
timestamp 1719641852
transform 1 0 2412 0 1 2905
box -2 -3 10 103
use OAI21X1  OAI21X1_644
timestamp 1719641852
transform 1 0 2420 0 1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_645
timestamp 1719641852
transform 1 0 2452 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_267
timestamp 1719641852
transform -1 0 2508 0 1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_601
timestamp 1719641852
transform -1 0 2540 0 1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_600
timestamp 1719641852
transform -1 0 2572 0 1 2905
box -2 -3 34 103
use DFFSR  DFFSR_166
timestamp 1719641852
transform -1 0 2748 0 1 2905
box -2 -3 178 103
use INVX2  INVX2_144
timestamp 1719641852
transform 1 0 2748 0 1 2905
box -2 -3 18 103
use DFFSR  DFFSR_196
timestamp 1719641852
transform -1 0 2940 0 1 2905
box -2 -3 178 103
use FILL  FILL_29_5_0
timestamp 1719641852
transform 1 0 2940 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_5_1
timestamp 1719641852
transform 1 0 2948 0 1 2905
box -2 -3 10 103
use DFFSR  DFFSR_247
timestamp 1719641852
transform 1 0 2956 0 1 2905
box -2 -3 178 103
use NAND2X1  NAND2X1_342
timestamp 1719641852
transform -1 0 3156 0 1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_151
timestamp 1719641852
transform -1 0 3180 0 1 2905
box -2 -3 26 103
use XNOR2X1  XNOR2X1_11
timestamp 1719641852
transform 1 0 3180 0 1 2905
box -2 -3 58 103
use AOI21X1  AOI21X1_33
timestamp 1719641852
transform -1 0 3268 0 1 2905
box -2 -3 34 103
use NAND3X1  NAND3X1_172
timestamp 1719641852
transform -1 0 3300 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_147
timestamp 1719641852
transform 1 0 3300 0 1 2905
box -2 -3 26 103
use NAND3X1  NAND3X1_187
timestamp 1719641852
transform -1 0 3356 0 1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_44
timestamp 1719641852
transform -1 0 3388 0 1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_277
timestamp 1719641852
transform 1 0 3388 0 1 2905
box -2 -3 34 103
use FILL  FILL_29_6_0
timestamp 1719641852
transform 1 0 3420 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_6_1
timestamp 1719641852
transform 1 0 3428 0 1 2905
box -2 -3 10 103
use NAND3X1  NAND3X1_190
timestamp 1719641852
transform 1 0 3436 0 1 2905
box -2 -3 34 103
use XNOR2X1  XNOR2X1_5
timestamp 1719641852
transform 1 0 3468 0 1 2905
box -2 -3 58 103
use NAND2X1  NAND2X1_128
timestamp 1719641852
transform 1 0 3524 0 1 2905
box -2 -3 26 103
use AND2X2  AND2X2_21
timestamp 1719641852
transform 1 0 3548 0 1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_32
timestamp 1719641852
transform 1 0 3580 0 1 2905
box -2 -3 34 103
use AOI22X1  AOI22X1_36
timestamp 1719641852
transform 1 0 3612 0 1 2905
box -2 -3 42 103
use NAND3X1  NAND3X1_198
timestamp 1719641852
transform 1 0 3652 0 1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_62
timestamp 1719641852
transform -1 0 3708 0 1 2905
box -2 -3 26 103
use AND2X2  AND2X2_11
timestamp 1719641852
transform -1 0 3740 0 1 2905
box -2 -3 34 103
use INVX1  INVX1_87
timestamp 1719641852
transform -1 0 3756 0 1 2905
box -2 -3 18 103
use NOR2X1  NOR2X1_67
timestamp 1719641852
transform 1 0 3756 0 1 2905
box -2 -3 26 103
use BUFX2  BUFX2_20
timestamp 1719641852
transform -1 0 28 0 -1 3105
box -2 -3 26 103
use DFFSR  DFFSR_64
timestamp 1719641852
transform -1 0 204 0 -1 3105
box -2 -3 178 103
use CLKBUF1  CLKBUF1_61
timestamp 1719641852
transform 1 0 4 0 1 3105
box -2 -3 74 103
use CLKBUF1  CLKBUF1_49
timestamp 1719641852
transform 1 0 76 0 1 3105
box -2 -3 74 103
use DFFSR  DFFSR_18
timestamp 1719641852
transform 1 0 148 0 1 3105
box -2 -3 178 103
use NOR2X1  NOR2X1_18
timestamp 1719641852
transform 1 0 204 0 -1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_144
timestamp 1719641852
transform 1 0 228 0 -1 3105
box -2 -3 34 103
use FILL  FILL_30_0_0
timestamp 1719641852
transform 1 0 260 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_0_1
timestamp 1719641852
transform 1 0 268 0 -1 3105
box -2 -3 10 103
use DFFSR  DFFSR_7
timestamp 1719641852
transform 1 0 276 0 -1 3105
box -2 -3 178 103
use FILL  FILL_31_0_0
timestamp 1719641852
transform 1 0 324 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_0_1
timestamp 1719641852
transform 1 0 332 0 1 3105
box -2 -3 10 103
use DFFSR  DFFSR_33
timestamp 1719641852
transform 1 0 340 0 1 3105
box -2 -3 178 103
use BUFX4  BUFX4_139
timestamp 1719641852
transform -1 0 484 0 -1 3105
box -2 -3 34 103
use INVX2  INVX2_15
timestamp 1719641852
transform 1 0 484 0 -1 3105
box -2 -3 18 103
use DFFSR  DFFSR_40
timestamp 1719641852
transform 1 0 500 0 -1 3105
box -2 -3 178 103
use DFFSR  DFFSR_1
timestamp 1719641852
transform 1 0 516 0 1 3105
box -2 -3 178 103
use OAI21X1  OAI21X1_62
timestamp 1719641852
transform -1 0 708 0 -1 3105
box -2 -3 34 103
use BUFX4  BUFX4_181
timestamp 1719641852
transform -1 0 740 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_50
timestamp 1719641852
transform 1 0 692 0 1 3105
box -2 -3 34 103
use NAND3X1  NAND3X1_27
timestamp 1719641852
transform -1 0 756 0 1 3105
box -2 -3 34 103
use NAND3X1  NAND3X1_28
timestamp 1719641852
transform 1 0 788 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_87
timestamp 1719641852
transform -1 0 788 0 1 3105
box -2 -3 34 103
use BUFX4  BUFX4_179
timestamp 1719641852
transform 1 0 804 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_51
timestamp 1719641852
transform 1 0 772 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_59
timestamp 1719641852
transform 1 0 740 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_26
timestamp 1719641852
transform 1 0 900 0 1 3105
box -2 -3 26 103
use NAND3X1  NAND3X1_12
timestamp 1719641852
transform 1 0 868 0 1 3105
box -2 -3 34 103
use FILL  FILL_31_1_1
timestamp 1719641852
transform 1 0 860 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_1_0
timestamp 1719641852
transform 1 0 852 0 1 3105
box -2 -3 10 103
use OAI21X1  OAI21X1_20
timestamp 1719641852
transform 1 0 820 0 1 3105
box -2 -3 34 103
use FILL  FILL_30_1_1
timestamp 1719641852
transform 1 0 876 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_1_0
timestamp 1719641852
transform 1 0 868 0 -1 3105
box -2 -3 10 103
use OAI21X1  OAI21X1_83
timestamp 1719641852
transform -1 0 868 0 -1 3105
box -2 -3 34 103
use DFFSR  DFFSR_35
timestamp 1719641852
transform 1 0 884 0 -1 3105
box -2 -3 178 103
use OAI21X1  OAI21X1_89
timestamp 1719641852
transform -1 0 1092 0 -1 3105
box -2 -3 34 103
use INVX1  INVX1_10
timestamp 1719641852
transform -1 0 940 0 1 3105
box -2 -3 18 103
use BUFX4  BUFX4_81
timestamp 1719641852
transform -1 0 972 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_19
timestamp 1719641852
transform 1 0 972 0 1 3105
box -2 -3 34 103
use DFFSR  DFFSR_38
timestamp 1719641852
transform 1 0 1004 0 1 3105
box -2 -3 178 103
use OAI21X1  OAI21X1_91
timestamp 1719641852
transform -1 0 1124 0 -1 3105
box -2 -3 34 103
use INVX1  INVX1_24
timestamp 1719641852
transform -1 0 1140 0 -1 3105
box -2 -3 18 103
use INVX2  INVX2_21
timestamp 1719641852
transform -1 0 1156 0 -1 3105
box -2 -3 18 103
use DFFSR  DFFSR_23
timestamp 1719641852
transform -1 0 1332 0 -1 3105
box -2 -3 178 103
use INVX2  INVX2_22
timestamp 1719641852
transform -1 0 1196 0 1 3105
box -2 -3 18 103
use DFFSR  DFFSR_21
timestamp 1719641852
transform 1 0 1196 0 1 3105
box -2 -3 178 103
use NAND2X1  NAND2X1_37
timestamp 1719641852
transform -1 0 1356 0 -1 3105
box -2 -3 26 103
use FILL  FILL_31_2_1
timestamp 1719641852
transform 1 0 1380 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_2_0
timestamp 1719641852
transform 1 0 1372 0 1 3105
box -2 -3 10 103
use NAND3X1  NAND3X1_74
timestamp 1719641852
transform 1 0 1372 0 -1 3105
box -2 -3 34 103
use FILL  FILL_30_2_1
timestamp 1719641852
transform 1 0 1364 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_2_0
timestamp 1719641852
transform 1 0 1356 0 -1 3105
box -2 -3 10 103
use OAI21X1  OAI21X1_26
timestamp 1719641852
transform 1 0 1404 0 1 3105
box -2 -3 34 103
use INVX1  INVX1_13
timestamp 1719641852
transform 1 0 1388 0 1 3105
box -2 -3 18 103
use NAND3X1  NAND3X1_70
timestamp 1719641852
transform 1 0 1404 0 -1 3105
box -2 -3 34 103
use NAND3X1  NAND3X1_15
timestamp 1719641852
transform 1 0 1436 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_30
timestamp 1719641852
transform 1 0 1436 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_13
timestamp 1719641852
transform 1 0 1524 0 1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_12
timestamp 1719641852
transform -1 0 1524 0 1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_25
timestamp 1719641852
transform 1 0 1468 0 1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_1
timestamp 1719641852
transform -1 0 1540 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_36
timestamp 1719641852
transform 1 0 1484 0 -1 3105
box -2 -3 26 103
use INVX1  INVX1_15
timestamp 1719641852
transform -1 0 1484 0 -1 3105
box -2 -3 18 103
use CLKBUF1  CLKBUF1_59
timestamp 1719641852
transform 1 0 1548 0 1 3105
box -2 -3 74 103
use NAND3X1  NAND3X1_91
timestamp 1719641852
transform 1 0 1604 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_29
timestamp 1719641852
transform 1 0 1572 0 -1 3105
box -2 -3 34 103
use NAND3X1  NAND3X1_17
timestamp 1719641852
transform 1 0 1540 0 -1 3105
box -2 -3 34 103
use BUFX4  BUFX4_161
timestamp 1719641852
transform -1 0 1652 0 1 3105
box -2 -3 34 103
use NAND3X1  NAND3X1_86
timestamp 1719641852
transform -1 0 1748 0 1 3105
box -2 -3 34 103
use BUFX4  BUFX4_165
timestamp 1719641852
transform -1 0 1716 0 1 3105
box -2 -3 34 103
use BUFX4  BUFX4_164
timestamp 1719641852
transform -1 0 1684 0 1 3105
box -2 -3 34 103
use AOI22X1  AOI22X1_2
timestamp 1719641852
transform 1 0 1692 0 -1 3105
box -2 -3 42 103
use NAND2X1  NAND2X1_65
timestamp 1719641852
transform -1 0 1692 0 -1 3105
box -2 -3 26 103
use BUFX4  BUFX4_134
timestamp 1719641852
transform 1 0 1636 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_10
timestamp 1719641852
transform 1 0 1796 0 1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_219
timestamp 1719641852
transform 1 0 1772 0 1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_60
timestamp 1719641852
transform -1 0 1772 0 1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_214
timestamp 1719641852
transform 1 0 1756 0 -1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_15
timestamp 1719641852
transform 1 0 1732 0 -1 3105
box -2 -3 26 103
use DFFSR  DFFSR_133
timestamp 1719641852
transform -1 0 1956 0 -1 3105
box -2 -3 178 103
use OAI21X1  OAI21X1_672
timestamp 1719641852
transform 1 0 1836 0 1 3105
box -2 -3 34 103
use INVX2  INVX2_161
timestamp 1719641852
transform 1 0 1820 0 1 3105
box -2 -3 18 103
use NAND2X1  NAND2X1_294
timestamp 1719641852
transform -1 0 1892 0 1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_673
timestamp 1719641852
transform -1 0 1940 0 1 3105
box -2 -3 34 103
use FILL  FILL_31_3_1
timestamp 1719641852
transform -1 0 1908 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_3_0
timestamp 1719641852
transform -1 0 1900 0 1 3105
box -2 -3 10 103
use NAND2X1  NAND2X1_293
timestamp 1719641852
transform 1 0 1940 0 1 3105
box -2 -3 26 103
use FILL  FILL_30_3_0
timestamp 1719641852
transform 1 0 1956 0 -1 3105
box -2 -3 10 103
use OAI21X1  OAI21X1_671
timestamp 1719641852
transform -1 0 1996 0 1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_264
timestamp 1719641852
transform 1 0 1972 0 -1 3105
box -2 -3 26 103
use FILL  FILL_30_3_1
timestamp 1719641852
transform 1 0 1964 0 -1 3105
box -2 -3 10 103
use OAI21X1  OAI21X1_589
timestamp 1719641852
transform -1 0 2052 0 1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_292
timestamp 1719641852
transform -1 0 2020 0 1 3105
box -2 -3 26 103
use INVX2  INVX2_54
timestamp 1719641852
transform 1 0 2020 0 -1 3105
box -2 -3 18 103
use NOR2X1  NOR2X1_308
timestamp 1719641852
transform -1 0 2020 0 -1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_226
timestamp 1719641852
transform 1 0 2052 0 1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_586
timestamp 1719641852
transform 1 0 2068 0 -1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_200
timestamp 1719641852
transform 1 0 2036 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_588
timestamp 1719641852
transform -1 0 2108 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_587
timestamp 1719641852
transform -1 0 2132 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_605
timestamp 1719641852
transform 1 0 2132 0 1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_317
timestamp 1719641852
transform -1 0 2132 0 1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_604
timestamp 1719641852
transform -1 0 2164 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_606
timestamp 1719641852
transform 1 0 2164 0 1 3105
box -2 -3 34 103
use INVX2  INVX2_147
timestamp 1719641852
transform 1 0 2164 0 -1 3105
box -2 -3 18 103
use OAI21X1  OAI21X1_650
timestamp 1719641852
transform -1 0 2228 0 1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_211
timestamp 1719641852
transform -1 0 2236 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_268
timestamp 1719641852
transform 1 0 2180 0 -1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_245
timestamp 1719641852
transform -1 0 2252 0 1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_603
timestamp 1719641852
transform -1 0 2268 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_651
timestamp 1719641852
transform -1 0 2308 0 1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_282
timestamp 1719641852
transform 1 0 2252 0 1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_649
timestamp 1719641852
transform -1 0 2300 0 -1 3105
box -2 -3 34 103
use INVX2  INVX2_100
timestamp 1719641852
transform 1 0 2308 0 1 3105
box -2 -3 18 103
use NOR2X1  NOR2X1_281
timestamp 1719641852
transform 1 0 2300 0 -1 3105
box -2 -3 26 103
use AOI21X1  AOI21X1_242
timestamp 1719641852
transform -1 0 2380 0 1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_304
timestamp 1719641852
transform 1 0 2324 0 1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_648
timestamp 1719641852
transform -1 0 2380 0 -1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_310
timestamp 1719641852
transform -1 0 2348 0 -1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_305
timestamp 1719641852
transform -1 0 2404 0 1 3105
box -2 -3 26 103
use NOR2X1  NOR2X1_312
timestamp 1719641852
transform 1 0 2380 0 -1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_690
timestamp 1719641852
transform -1 0 2452 0 1 3105
box -2 -3 34 103
use FILL  FILL_31_4_1
timestamp 1719641852
transform -1 0 2420 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_4_0
timestamp 1719641852
transform -1 0 2412 0 1 3105
box -2 -3 10 103
use NOR2X1  NOR2X1_282
timestamp 1719641852
transform 1 0 2420 0 -1 3105
box -2 -3 26 103
use FILL  FILL_30_4_1
timestamp 1719641852
transform 1 0 2412 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_4_0
timestamp 1719641852
transform 1 0 2404 0 -1 3105
box -2 -3 10 103
use INVX2  INVX2_107
timestamp 1719641852
transform 1 0 2452 0 1 3105
box -2 -3 18 103
use OAI21X1  OAI21X1_732
timestamp 1719641852
transform -1 0 2476 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_716
timestamp 1719641852
transform 1 0 2484 0 1 3105
box -2 -3 34 103
use INVX1  INVX1_158
timestamp 1719641852
transform 1 0 2468 0 1 3105
box -2 -3 18 103
use OAI21X1  OAI21X1_646
timestamp 1719641852
transform 1 0 2500 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_326
timestamp 1719641852
transform -1 0 2500 0 -1 3105
box -2 -3 26 103
use NOR2X1  NOR2X1_320
timestamp 1719641852
transform 1 0 2516 0 1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_647
timestamp 1719641852
transform 1 0 2532 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_609
timestamp 1719641852
transform -1 0 2636 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_610
timestamp 1719641852
transform -1 0 2604 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_717
timestamp 1719641852
transform 1 0 2540 0 1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_212
timestamp 1719641852
transform 1 0 2612 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_316
timestamp 1719641852
transform 1 0 2588 0 -1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_281
timestamp 1719641852
transform -1 0 2588 0 -1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_269
timestamp 1719641852
transform -1 0 2692 0 1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_611
timestamp 1719641852
transform 1 0 2636 0 1 3105
box -2 -3 34 103
use INVX2  INVX2_103
timestamp 1719641852
transform 1 0 2700 0 -1 3105
box -2 -3 18 103
use NAND2X1  NAND2X1_324
timestamp 1719641852
transform 1 0 2676 0 -1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_608
timestamp 1719641852
transform -1 0 2676 0 -1 3105
box -2 -3 34 103
use DFFSR  DFFSR_121
timestamp 1719641852
transform 1 0 2692 0 1 3105
box -2 -3 178 103
use DFFSR  DFFSR_149
timestamp 1719641852
transform -1 0 2892 0 -1 3105
box -2 -3 178 103
use FILL  FILL_30_5_0
timestamp 1719641852
transform -1 0 2900 0 -1 3105
box -2 -3 10 103
use BUFX4  BUFX4_109
timestamp 1719641852
transform -1 0 2900 0 1 3105
box -2 -3 34 103
use XNOR2X1  XNOR2X1_4
timestamp 1719641852
transform 1 0 2940 0 1 3105
box -2 -3 58 103
use INVX4  INVX4_2
timestamp 1719641852
transform -1 0 2940 0 1 3105
box -2 -3 26 103
use FILL  FILL_31_5_1
timestamp 1719641852
transform -1 0 2916 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_5_0
timestamp 1719641852
transform -1 0 2908 0 1 3105
box -2 -3 10 103
use CLKBUF1  CLKBUF1_6
timestamp 1719641852
transform -1 0 2980 0 -1 3105
box -2 -3 74 103
use FILL  FILL_30_5_1
timestamp 1719641852
transform -1 0 2908 0 -1 3105
box -2 -3 10 103
use XNOR2X1  XNOR2X1_10
timestamp 1719641852
transform 1 0 3020 0 1 3105
box -2 -3 58 103
use NAND2X1  NAND2X1_132
timestamp 1719641852
transform 1 0 2996 0 1 3105
box -2 -3 26 103
use OAI22X1  OAI22X1_42
timestamp 1719641852
transform 1 0 3052 0 -1 3105
box -2 -3 42 103
use CLKBUF1  CLKBUF1_48
timestamp 1719641852
transform 1 0 2980 0 -1 3105
box -2 -3 74 103
use AOI21X1  AOI21X1_47
timestamp 1719641852
transform 1 0 3076 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_282
timestamp 1719641852
transform -1 0 3140 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_792
timestamp 1719641852
transform -1 0 3124 0 -1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_48
timestamp 1719641852
transform 1 0 3140 0 1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_150
timestamp 1719641852
transform -1 0 3164 0 -1 3105
box -2 -3 26 103
use INVX2  INVX2_46
timestamp 1719641852
transform -1 0 3140 0 -1 3105
box -2 -3 18 103
use OAI21X1  OAI21X1_281
timestamp 1719641852
transform -1 0 3204 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_280
timestamp 1719641852
transform -1 0 3196 0 -1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_47
timestamp 1719641852
transform -1 0 3252 0 1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_136
timestamp 1719641852
transform 1 0 3204 0 1 3105
box -2 -3 26 103
use NOR2X1  NOR2X1_340
timestamp 1719641852
transform 1 0 3212 0 -1 3105
box -2 -3 26 103
use INVX1  INVX1_107
timestamp 1719641852
transform -1 0 3212 0 -1 3105
box -2 -3 18 103
use OAI21X1  OAI21X1_273
timestamp 1719641852
transform 1 0 3252 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_269
timestamp 1719641852
transform -1 0 3268 0 -1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_55
timestamp 1719641852
transform 1 0 3284 0 1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_190
timestamp 1719641852
transform 1 0 3268 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_105
timestamp 1719641852
transform 1 0 3324 0 1 3105
box -2 -3 26 103
use INVX1  INVX1_85
timestamp 1719641852
transform -1 0 3324 0 1 3105
box -2 -3 18 103
use NOR2X1  NOR2X1_53
timestamp 1719641852
transform -1 0 3356 0 -1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_189
timestamp 1719641852
transform 1 0 3300 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_192
timestamp 1719641852
transform -1 0 3380 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_188
timestamp 1719641852
transform 1 0 3372 0 -1 3105
box -2 -3 34 103
use INVX2  INVX2_45
timestamp 1719641852
transform 1 0 3356 0 -1 3105
box -2 -3 18 103
use NAND2X1  NAND2X1_148
timestamp 1719641852
transform 1 0 3396 0 1 3105
box -2 -3 26 103
use INVX1  INVX1_108
timestamp 1719641852
transform -1 0 3396 0 1 3105
box -2 -3 18 103
use FILL  FILL_30_6_0
timestamp 1719641852
transform 1 0 3404 0 -1 3105
box -2 -3 10 103
use AND2X2  AND2X2_10
timestamp 1719641852
transform 1 0 3436 0 1 3105
box -2 -3 34 103
use FILL  FILL_31_6_1
timestamp 1719641852
transform 1 0 3428 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_6_0
timestamp 1719641852
transform 1 0 3420 0 1 3105
box -2 -3 10 103
use OAI21X1  OAI21X1_194
timestamp 1719641852
transform 1 0 3420 0 -1 3105
box -2 -3 34 103
use FILL  FILL_30_6_1
timestamp 1719641852
transform 1 0 3412 0 -1 3105
box -2 -3 10 103
use NOR2X1  NOR2X1_58
timestamp 1719641852
transform -1 0 3492 0 1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_193
timestamp 1719641852
transform 1 0 3452 0 -1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_28
timestamp 1719641852
transform 1 0 3508 0 1 3105
box -2 -3 34 103
use INVX1  INVX1_88
timestamp 1719641852
transform -1 0 3508 0 1 3105
box -2 -3 18 103
use OAI21X1  OAI21X1_276
timestamp 1719641852
transform 1 0 3508 0 -1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_59
timestamp 1719641852
transform 1 0 3484 0 -1 3105
box -2 -3 26 103
use NAND3X1  NAND3X1_184
timestamp 1719641852
transform -1 0 3572 0 1 3105
box -2 -3 34 103
use NAND3X1  NAND3X1_193
timestamp 1719641852
transform -1 0 3572 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_146
timestamp 1719641852
transform 1 0 3572 0 1 3105
box -2 -3 26 103
use NAND3X1  NAND3X1_191
timestamp 1719641852
transform -1 0 3604 0 -1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_51
timestamp 1719641852
transform 1 0 3620 0 1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_153
timestamp 1719641852
transform 1 0 3596 0 1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_288
timestamp 1719641852
transform -1 0 3636 0 -1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_54
timestamp 1719641852
transform 1 0 3652 0 1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_41
timestamp 1719641852
transform -1 0 3668 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_144
timestamp 1719641852
transform 1 0 3684 0 1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_292
timestamp 1719641852
transform 1 0 3668 0 -1 3105
box -2 -3 34 103
use NAND3X1  NAND3X1_182
timestamp 1719641852
transform 1 0 3708 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_275
timestamp 1719641852
transform 1 0 3716 0 -1 3105
box -2 -3 34 103
use INVX1  INVX1_105
timestamp 1719641852
transform -1 0 3716 0 -1 3105
box -2 -3 18 103
use FILL  FILL_32_2
timestamp 1719641852
transform 1 0 3764 0 1 3105
box -2 -3 10 103
use FILL  FILL_32_1
timestamp 1719641852
transform 1 0 3756 0 1 3105
box -2 -3 10 103
use INVX1  INVX1_116
timestamp 1719641852
transform -1 0 3756 0 1 3105
box -2 -3 18 103
use NOR2X1  NOR2X1_66
timestamp 1719641852
transform -1 0 3772 0 -1 3105
box -2 -3 26 103
use FILL  FILL_32_3
timestamp 1719641852
transform 1 0 3772 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_1
timestamp 1719641852
transform -1 0 3780 0 -1 3105
box -2 -3 10 103
use BUFX2  BUFX2_37
timestamp 1719641852
transform -1 0 28 0 -1 3305
box -2 -3 26 103
use DFFSR  DFFSR_66
timestamp 1719641852
transform -1 0 204 0 -1 3305
box -2 -3 178 103
use BUFX4  BUFX4_93
timestamp 1719641852
transform 1 0 204 0 -1 3305
box -2 -3 34 103
use DFFSR  DFFSR_6
timestamp 1719641852
transform 1 0 236 0 -1 3305
box -2 -3 178 103
use FILL  FILL_32_0_0
timestamp 1719641852
transform -1 0 420 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_0_1
timestamp 1719641852
transform -1 0 428 0 -1 3305
box -2 -3 10 103
use NAND2X1  NAND2X1_77
timestamp 1719641852
transform -1 0 452 0 -1 3305
box -2 -3 26 103
use OAI21X1  OAI21X1_133
timestamp 1719641852
transform -1 0 484 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_131
timestamp 1719641852
transform 1 0 484 0 -1 3305
box -2 -3 34 103
use INVX2  INVX2_14
timestamp 1719641852
transform 1 0 516 0 -1 3305
box -2 -3 18 103
use INVX1  INVX1_21
timestamp 1719641852
transform 1 0 532 0 -1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_76
timestamp 1719641852
transform 1 0 548 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_77
timestamp 1719641852
transform 1 0 580 0 -1 3305
box -2 -3 34 103
use INVX2  INVX2_11
timestamp 1719641852
transform 1 0 612 0 -1 3305
box -2 -3 18 103
use BUFX4  BUFX4_92
timestamp 1719641852
transform 1 0 628 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_54
timestamp 1719641852
transform -1 0 692 0 -1 3305
box -2 -3 34 103
use INVX2  INVX2_9
timestamp 1719641852
transform 1 0 692 0 -1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_60
timestamp 1719641852
transform 1 0 708 0 -1 3305
box -2 -3 34 103
use NAND3X1  NAND3X1_32
timestamp 1719641852
transform -1 0 772 0 -1 3305
box -2 -3 34 103
use INVX2  INVX2_10
timestamp 1719641852
transform 1 0 772 0 -1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_52
timestamp 1719641852
transform -1 0 820 0 -1 3305
box -2 -3 34 103
use INVX2  INVX2_20
timestamp 1719641852
transform -1 0 836 0 -1 3305
box -2 -3 18 103
use FILL  FILL_32_1_0
timestamp 1719641852
transform -1 0 844 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_1_1
timestamp 1719641852
transform -1 0 852 0 -1 3305
box -2 -3 10 103
use DFFSR  DFFSR_24
timestamp 1719641852
transform -1 0 1028 0 -1 3305
box -2 -3 178 103
use DFFSR  DFFSR_39
timestamp 1719641852
transform 1 0 1028 0 -1 3305
box -2 -3 178 103
use OAI21X1  OAI21X1_28
timestamp 1719641852
transform 1 0 1204 0 -1 3305
box -2 -3 34 103
use INVX1  INVX1_14
timestamp 1719641852
transform 1 0 1236 0 -1 3305
box -2 -3 18 103
use NAND3X1  NAND3X1_16
timestamp 1719641852
transform 1 0 1252 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_27
timestamp 1719641852
transform 1 0 1284 0 -1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_14
timestamp 1719641852
transform 1 0 1316 0 -1 3305
box -2 -3 26 103
use OAI21X1  OAI21X1_145
timestamp 1719641852
transform 1 0 1340 0 -1 3305
box -2 -3 34 103
use FILL  FILL_32_2_0
timestamp 1719641852
transform -1 0 1380 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_2_1
timestamp 1719641852
transform -1 0 1388 0 -1 3305
box -2 -3 10 103
use NAND3X1  NAND3X1_14
timestamp 1719641852
transform -1 0 1420 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_24
timestamp 1719641852
transform -1 0 1452 0 -1 3305
box -2 -3 34 103
use INVX1  INVX1_12
timestamp 1719641852
transform -1 0 1468 0 -1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_23
timestamp 1719641852
transform 1 0 1468 0 -1 3305
box -2 -3 34 103
use BUFX4  BUFX4_100
timestamp 1719641852
transform -1 0 1532 0 -1 3305
box -2 -3 34 103
use CLKBUF1  CLKBUF1_44
timestamp 1719641852
transform -1 0 1604 0 -1 3305
box -2 -3 74 103
use BUFX4  BUFX4_160
timestamp 1719641852
transform -1 0 1636 0 -1 3305
box -2 -3 34 103
use BUFX4  BUFX4_162
timestamp 1719641852
transform -1 0 1668 0 -1 3305
box -2 -3 34 103
use BUFX4  BUFX4_163
timestamp 1719641852
transform -1 0 1700 0 -1 3305
box -2 -3 34 103
use DFFSR  DFFSR_137
timestamp 1719641852
transform -1 0 1876 0 -1 3305
box -2 -3 178 103
use FILL  FILL_32_3_0
timestamp 1719641852
transform -1 0 1884 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_3_1
timestamp 1719641852
transform -1 0 1892 0 -1 3305
box -2 -3 10 103
use NAND2X1  NAND2X1_216
timestamp 1719641852
transform -1 0 1916 0 -1 3305
box -2 -3 26 103
use DFFSR  DFFSR_170
timestamp 1719641852
transform -1 0 2092 0 -1 3305
box -2 -3 178 103
use DFFSR  DFFSR_165
timestamp 1719641852
transform -1 0 2268 0 -1 3305
box -2 -3 178 103
use OAI21X1  OAI21X1_691
timestamp 1719641852
transform -1 0 2300 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_692
timestamp 1719641852
transform 1 0 2300 0 -1 3305
box -2 -3 34 103
use INVX1  INVX1_153
timestamp 1719641852
transform -1 0 2348 0 -1 3305
box -2 -3 18 103
use NOR2X1  NOR2X1_313
timestamp 1719641852
transform 1 0 2348 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_327
timestamp 1719641852
transform 1 0 2372 0 -1 3305
box -2 -3 26 103
use FILL  FILL_32_4_0
timestamp 1719641852
transform 1 0 2396 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_4_1
timestamp 1719641852
transform 1 0 2404 0 -1 3305
box -2 -3 10 103
use OAI21X1  OAI21X1_733
timestamp 1719641852
transform 1 0 2412 0 -1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_324
timestamp 1719641852
transform 1 0 2444 0 -1 3305
box -2 -3 26 103
use OAI21X1  OAI21X1_734
timestamp 1719641852
transform 1 0 2468 0 -1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_325
timestamp 1719641852
transform -1 0 2524 0 -1 3305
box -2 -3 26 103
use INVX1  INVX1_160
timestamp 1719641852
transform 1 0 2524 0 -1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_730
timestamp 1719641852
transform 1 0 2540 0 -1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_323
timestamp 1719641852
transform 1 0 2572 0 -1 3305
box -2 -3 26 103
use OAI21X1  OAI21X1_731
timestamp 1719641852
transform 1 0 2596 0 -1 3305
box -2 -3 34 103
use BUFX4  BUFX4_130
timestamp 1719641852
transform -1 0 2660 0 -1 3305
box -2 -3 34 103
use BUFX4  BUFX4_132
timestamp 1719641852
transform 1 0 2660 0 -1 3305
box -2 -3 34 103
use DFFSR  DFFSR_164
timestamp 1719641852
transform -1 0 2868 0 -1 3305
box -2 -3 178 103
use XOR2X1  XOR2X1_3
timestamp 1719641852
transform -1 0 2924 0 -1 3305
box -2 -3 58 103
use FILL  FILL_32_5_0
timestamp 1719641852
transform -1 0 2932 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_5_1
timestamp 1719641852
transform -1 0 2940 0 -1 3305
box -2 -3 10 103
use INVX4  INVX4_11
timestamp 1719641852
transform -1 0 2964 0 -1 3305
box -2 -3 26 103
use INVX4  INVX4_3
timestamp 1719641852
transform 1 0 2964 0 -1 3305
box -2 -3 26 103
use NOR2X1  NOR2X1_342
timestamp 1719641852
transform -1 0 3012 0 -1 3305
box -2 -3 26 103
use OAI21X1  OAI21X1_793
timestamp 1719641852
transform -1 0 3044 0 -1 3305
box -2 -3 34 103
use INVX2  INVX2_53
timestamp 1719641852
transform 1 0 3044 0 -1 3305
box -2 -3 18 103
use BUFX4  BUFX4_112
timestamp 1719641852
transform 1 0 3060 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_187
timestamp 1719641852
transform -1 0 3124 0 -1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_104
timestamp 1719641852
transform 1 0 3124 0 -1 3305
box -2 -3 26 103
use OAI21X1  OAI21X1_283
timestamp 1719641852
transform 1 0 3148 0 -1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_101
timestamp 1719641852
transform 1 0 3180 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_135
timestamp 1719641852
transform 1 0 3204 0 -1 3305
box -2 -3 26 103
use OAI21X1  OAI21X1_271
timestamp 1719641852
transform 1 0 3228 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_270
timestamp 1719641852
transform -1 0 3292 0 -1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_175
timestamp 1719641852
transform -1 0 3316 0 -1 3305
box -2 -3 26 103
use AND2X2  AND2X2_9
timestamp 1719641852
transform -1 0 3348 0 -1 3305
box -2 -3 34 103
use AOI21X1  AOI21X1_35
timestamp 1719641852
transform -1 0 3380 0 -1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_137
timestamp 1719641852
transform -1 0 3404 0 -1 3305
box -2 -3 26 103
use FILL  FILL_32_6_0
timestamp 1719641852
transform 1 0 3404 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_6_1
timestamp 1719641852
transform 1 0 3412 0 -1 3305
box -2 -3 10 103
use NAND3X1  NAND3X1_188
timestamp 1719641852
transform 1 0 3420 0 -1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_57
timestamp 1719641852
transform -1 0 3476 0 -1 3305
box -2 -3 26 103
use NOR2X1  NOR2X1_56
timestamp 1719641852
transform 1 0 3476 0 -1 3305
box -2 -3 26 103
use AOI21X1  AOI21X1_53
timestamp 1719641852
transform -1 0 3532 0 -1 3305
box -2 -3 34 103
use NAND3X1  NAND3X1_197
timestamp 1719641852
transform 1 0 3532 0 -1 3305
box -2 -3 34 103
use NAND3X1  NAND3X1_185
timestamp 1719641852
transform -1 0 3596 0 -1 3305
box -2 -3 34 103
use NAND3X1  NAND3X1_192
timestamp 1719641852
transform -1 0 3628 0 -1 3305
box -2 -3 34 103
use AOI21X1  AOI21X1_45
timestamp 1719641852
transform -1 0 3660 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_278
timestamp 1719641852
transform -1 0 3692 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_290
timestamp 1719641852
transform 1 0 3692 0 -1 3305
box -2 -3 34 103
use AOI21X1  AOI21X1_39
timestamp 1719641852
transform 1 0 3724 0 -1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_179
timestamp 1719641852
transform 1 0 3756 0 -1 3305
box -2 -3 26 103
use BUFX2  BUFX2_35
timestamp 1719641852
transform -1 0 28 0 1 3305
box -2 -3 26 103
use BUFX2  BUFX2_69
timestamp 1719641852
transform -1 0 52 0 1 3305
box -2 -3 26 103
use INVX1  INVX1_64
timestamp 1719641852
transform 1 0 52 0 1 3305
box -2 -3 18 103
use DFFSR  DFFSR_63
timestamp 1719641852
transform -1 0 244 0 1 3305
box -2 -3 178 103
use OAI22X1  OAI22X1_39
timestamp 1719641852
transform 1 0 244 0 1 3305
box -2 -3 42 103
use OAI21X1  OAI21X1_132
timestamp 1719641852
transform 1 0 284 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_150
timestamp 1719641852
transform 1 0 316 0 1 3305
box -2 -3 34 103
use FILL  FILL_33_0_0
timestamp 1719641852
transform 1 0 348 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_0_1
timestamp 1719641852
transform 1 0 356 0 1 3305
box -2 -3 10 103
use OAI21X1  OAI21X1_129
timestamp 1719641852
transform 1 0 364 0 1 3305
box -2 -3 34 103
use BUFX4  BUFX4_144
timestamp 1719641852
transform -1 0 428 0 1 3305
box -2 -3 34 103
use DFFSR  DFFSR_3
timestamp 1719641852
transform -1 0 604 0 1 3305
box -2 -3 178 103
use NAND2X1  NAND2X1_33
timestamp 1719641852
transform -1 0 628 0 1 3305
box -2 -3 26 103
use OAI21X1  OAI21X1_127
timestamp 1719641852
transform -1 0 660 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_128
timestamp 1719641852
transform 1 0 660 0 1 3305
box -2 -3 34 103
use DFFSR  DFFSR_2
timestamp 1719641852
transform -1 0 868 0 1 3305
box -2 -3 178 103
use FILL  FILL_33_1_0
timestamp 1719641852
transform 1 0 868 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_1_1
timestamp 1719641852
transform 1 0 876 0 1 3305
box -2 -3 10 103
use BUFX4  BUFX4_145
timestamp 1719641852
transform 1 0 884 0 1 3305
box -2 -3 34 103
use NAND3X1  NAND3X1_18
timestamp 1719641852
transform -1 0 948 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_32
timestamp 1719641852
transform -1 0 980 0 1 3305
box -2 -3 34 103
use INVX1  INVX1_16
timestamp 1719641852
transform 1 0 980 0 1 3305
box -2 -3 18 103
use BUFX4  BUFX4_146
timestamp 1719641852
transform 1 0 996 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_31
timestamp 1719641852
transform 1 0 1028 0 1 3305
box -2 -3 34 103
use BUFX2  BUFX2_39
timestamp 1719641852
transform -1 0 1084 0 1 3305
box -2 -3 26 103
use DFFSR  DFFSR_81
timestamp 1719641852
transform -1 0 1260 0 1 3305
box -2 -3 178 103
use OAI21X1  OAI21X1_18
timestamp 1719641852
transform 1 0 1260 0 1 3305
box -2 -3 34 103
use NAND3X1  NAND3X1_11
timestamp 1719641852
transform 1 0 1292 0 1 3305
box -2 -3 34 103
use INVX1  INVX1_9
timestamp 1719641852
transform 1 0 1324 0 1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_17
timestamp 1719641852
transform 1 0 1340 0 1 3305
box -2 -3 34 103
use FILL  FILL_33_2_0
timestamp 1719641852
transform -1 0 1380 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_2_1
timestamp 1719641852
transform -1 0 1388 0 1 3305
box -2 -3 10 103
use DFFSR  DFFSR_20
timestamp 1719641852
transform -1 0 1564 0 1 3305
box -2 -3 178 103
use BUFX2  BUFX2_21
timestamp 1719641852
transform 1 0 1564 0 1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_16
timestamp 1719641852
transform 1 0 1588 0 1 3305
box -2 -3 26 103
use CLKBUF1  CLKBUF1_4
timestamp 1719641852
transform -1 0 1684 0 1 3305
box -2 -3 74 103
use CLKBUF1  CLKBUF1_29
timestamp 1719641852
transform 1 0 1684 0 1 3305
box -2 -3 74 103
use BUFX4  BUFX4_159
timestamp 1719641852
transform 1 0 1756 0 1 3305
box -2 -3 34 103
use DFFSR  DFFSR_83
timestamp 1719641852
transform 1 0 1788 0 1 3305
box -2 -3 178 103
use FILL  FILL_33_3_0
timestamp 1719641852
transform -1 0 1972 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_3_1
timestamp 1719641852
transform -1 0 1980 0 1 3305
box -2 -3 10 103
use NAND2X1  NAND2X1_9
timestamp 1719641852
transform -1 0 2004 0 1 3305
box -2 -3 26 103
use DFFSR  DFFSR_180
timestamp 1719641852
transform -1 0 2180 0 1 3305
box -2 -3 178 103
use NOR2X1  NOR2X1_348
timestamp 1719641852
transform -1 0 2204 0 1 3305
box -2 -3 26 103
use DFFSR  DFFSR_148
timestamp 1719641852
transform -1 0 2380 0 1 3305
box -2 -3 178 103
use NAND2X1  NAND2X1_229
timestamp 1719641852
transform 1 0 2380 0 1 3305
box -2 -3 26 103
use FILL  FILL_33_4_0
timestamp 1719641852
transform -1 0 2412 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_4_1
timestamp 1719641852
transform -1 0 2420 0 1 3305
box -2 -3 10 103
use INVX1  INVX1_161
timestamp 1719641852
transform -1 0 2436 0 1 3305
box -2 -3 18 103
use DFFSR  DFFSR_116
timestamp 1719641852
transform -1 0 2612 0 1 3305
box -2 -3 178 103
use DFFSR  DFFSR_248
timestamp 1719641852
transform 1 0 2612 0 1 3305
box -2 -3 178 103
use CLKBUF1  CLKBUF1_65
timestamp 1719641852
transform 1 0 2788 0 1 3305
box -2 -3 74 103
use OAI22X1  OAI22X1_43
timestamp 1719641852
transform 1 0 2860 0 1 3305
box -2 -3 42 103
use FILL  FILL_33_5_0
timestamp 1719641852
transform -1 0 2908 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_5_1
timestamp 1719641852
transform -1 0 2916 0 1 3305
box -2 -3 10 103
use NOR2X1  NOR2X1_341
timestamp 1719641852
transform -1 0 2940 0 1 3305
box -2 -3 26 103
use OAI22X1  OAI22X1_45
timestamp 1719641852
transform 1 0 2940 0 1 3305
box -2 -3 42 103
use NOR2X1  NOR2X1_343
timestamp 1719641852
transform 1 0 2980 0 1 3305
box -2 -3 26 103
use OAI21X1  OAI21X1_797
timestamp 1719641852
transform -1 0 3036 0 1 3305
box -2 -3 34 103
use XNOR2X1  XNOR2X1_8
timestamp 1719641852
transform 1 0 3036 0 1 3305
box -2 -3 58 103
use NAND3X1  NAND3X1_173
timestamp 1719641852
transform -1 0 3124 0 1 3305
box -2 -3 34 103
use OR2X2  OR2X2_8
timestamp 1719641852
transform -1 0 3156 0 1 3305
box -2 -3 34 103
use INVX2  INVX2_43
timestamp 1719641852
transform -1 0 3172 0 1 3305
box -2 -3 18 103
use NAND2X1  NAND2X1_134
timestamp 1719641852
transform -1 0 3196 0 1 3305
box -2 -3 26 103
use NAND3X1  NAND3X1_186
timestamp 1719641852
transform -1 0 3228 0 1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_133
timestamp 1719641852
transform 1 0 3228 0 1 3305
box -2 -3 26 103
use NAND3X1  NAND3X1_170
timestamp 1719641852
transform -1 0 3284 0 1 3305
box -2 -3 34 103
use INVX1  INVX1_103
timestamp 1719641852
transform -1 0 3300 0 1 3305
box -2 -3 18 103
use NAND3X1  NAND3X1_171
timestamp 1719641852
transform -1 0 3332 0 1 3305
box -2 -3 34 103
use INVX2  INVX2_48
timestamp 1719641852
transform -1 0 3348 0 1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_268
timestamp 1719641852
transform 1 0 3348 0 1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_272
timestamp 1719641852
transform 1 0 3380 0 1 3305
box -2 -3 34 103
use FILL  FILL_33_6_0
timestamp 1719641852
transform 1 0 3412 0 1 3305
box -2 -3 10 103
use FILL  FILL_33_6_1
timestamp 1719641852
transform 1 0 3420 0 1 3305
box -2 -3 10 103
use NAND3X1  NAND3X1_189
timestamp 1719641852
transform 1 0 3428 0 1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_129
timestamp 1719641852
transform 1 0 3460 0 1 3305
box -2 -3 26 103
use NOR2X1  NOR2X1_180
timestamp 1719641852
transform -1 0 3508 0 1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_130
timestamp 1719641852
transform 1 0 3508 0 1 3305
box -2 -3 26 103
use AOI21X1  AOI21X1_43
timestamp 1719641852
transform -1 0 3564 0 1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_145
timestamp 1719641852
transform -1 0 3588 0 1 3305
box -2 -3 26 103
use AND2X2  AND2X2_20
timestamp 1719641852
transform 1 0 3588 0 1 3305
box -2 -3 34 103
use AOI21X1  AOI21X1_37
timestamp 1719641852
transform 1 0 3620 0 1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_65
timestamp 1719641852
transform 1 0 3652 0 1 3305
box -2 -3 26 103
use AOI21X1  AOI21X1_38
timestamp 1719641852
transform 1 0 3676 0 1 3305
box -2 -3 34 103
use INVX2  INVX2_50
timestamp 1719641852
transform -1 0 3724 0 1 3305
box -2 -3 18 103
use NAND2X1  NAND2X1_141
timestamp 1719641852
transform -1 0 3748 0 1 3305
box -2 -3 26 103
use NAND3X1  NAND3X1_177
timestamp 1719641852
transform 1 0 3748 0 1 3305
box -2 -3 34 103
use BUFX2  BUFX2_26
timestamp 1719641852
transform -1 0 28 0 -1 3505
box -2 -3 26 103
use CLKBUF1  CLKBUF1_37
timestamp 1719641852
transform 1 0 28 0 -1 3505
box -2 -3 74 103
use CLKBUF1  CLKBUF1_15
timestamp 1719641852
transform 1 0 100 0 -1 3505
box -2 -3 74 103
use BUFX4  BUFX4_103
timestamp 1719641852
transform -1 0 204 0 -1 3505
box -2 -3 34 103
use BUFX2  BUFX2_48
timestamp 1719641852
transform -1 0 228 0 -1 3505
box -2 -3 26 103
use DFFSR  DFFSR_77
timestamp 1719641852
transform -1 0 404 0 -1 3505
box -2 -3 178 103
use FILL  FILL_34_0_0
timestamp 1719641852
transform -1 0 412 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_0_1
timestamp 1719641852
transform -1 0 420 0 -1 3505
box -2 -3 10 103
use BUFX2  BUFX2_3
timestamp 1719641852
transform -1 0 444 0 -1 3505
box -2 -3 26 103
use DFFSR  DFFSR_41
timestamp 1719641852
transform -1 0 620 0 -1 3505
box -2 -3 178 103
use DFFSR  DFFSR_37
timestamp 1719641852
transform 1 0 620 0 -1 3505
box -2 -3 178 103
use FILL  FILL_34_1_0
timestamp 1719641852
transform 1 0 796 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_1_1
timestamp 1719641852
transform 1 0 804 0 -1 3505
box -2 -3 10 103
use DFFSR  DFFSR_22
timestamp 1719641852
transform 1 0 812 0 -1 3505
box -2 -3 178 103
use DFFSR  DFFSR_17
timestamp 1719641852
transform 1 0 988 0 -1 3505
box -2 -3 178 103
use BUFX2  BUFX2_19
timestamp 1719641852
transform -1 0 1188 0 -1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_143
timestamp 1719641852
transform -1 0 1220 0 -1 3505
box -2 -3 34 103
use NOR2X1  NOR2X1_350
timestamp 1719641852
transform -1 0 1244 0 -1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_148
timestamp 1719641852
transform 1 0 1244 0 -1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_146
timestamp 1719641852
transform 1 0 1276 0 -1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_147
timestamp 1719641852
transform 1 0 1308 0 -1 3505
box -2 -3 34 103
use FILL  FILL_34_2_0
timestamp 1719641852
transform 1 0 1340 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_2_1
timestamp 1719641852
transform 1 0 1348 0 -1 3505
box -2 -3 10 103
use DFFSR  DFFSR_42
timestamp 1719641852
transform 1 0 1356 0 -1 3505
box -2 -3 178 103
use DFFSR  DFFSR_86
timestamp 1719641852
transform 1 0 1532 0 -1 3505
box -2 -3 178 103
use DFFSR  DFFSR_245
timestamp 1719641852
transform -1 0 1884 0 -1 3505
box -2 -3 178 103
use FILL  FILL_34_3_0
timestamp 1719641852
transform -1 0 1892 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_3_1
timestamp 1719641852
transform -1 0 1900 0 -1 3505
box -2 -3 10 103
use DFFSR  DFFSR_132
timestamp 1719641852
transform -1 0 2076 0 -1 3505
box -2 -3 178 103
use CLKBUF1  CLKBUF1_22
timestamp 1719641852
transform -1 0 2148 0 -1 3505
box -2 -3 74 103
use BUFX4  BUFX4_101
timestamp 1719641852
transform 1 0 2148 0 -1 3505
box -2 -3 34 103
use NOR2X1  NOR2X1_344
timestamp 1719641852
transform 1 0 2180 0 -1 3505
box -2 -3 26 103
use AND2X2  AND2X2_33
timestamp 1719641852
transform 1 0 2204 0 -1 3505
box -2 -3 34 103
use AOI21X1  AOI21X1_268
timestamp 1719641852
transform -1 0 2268 0 -1 3505
box -2 -3 34 103
use NOR2X1  NOR2X1_345
timestamp 1719641852
transform 1 0 2268 0 -1 3505
box -2 -3 26 103
use INVX1  INVX1_79
timestamp 1719641852
transform -1 0 2308 0 -1 3505
box -2 -3 18 103
use NOR2X1  NOR2X1_50
timestamp 1719641852
transform -1 0 2332 0 -1 3505
box -2 -3 26 103
use FILL  FILL_34_4_0
timestamp 1719641852
transform -1 0 2340 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_4_1
timestamp 1719641852
transform -1 0 2348 0 -1 3505
box -2 -3 10 103
use DFFSR  DFFSR_117
timestamp 1719641852
transform -1 0 2524 0 -1 3505
box -2 -3 178 103
use NOR2X1  NOR2X1_49
timestamp 1719641852
transform 1 0 2524 0 -1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_798
timestamp 1719641852
transform -1 0 2580 0 -1 3505
box -2 -3 34 103
use DFFSR  DFFSR_251
timestamp 1719641852
transform 1 0 2580 0 -1 3505
box -2 -3 178 103
use BUFX4  BUFX4_111
timestamp 1719641852
transform 1 0 2756 0 -1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_794
timestamp 1719641852
transform 1 0 2788 0 -1 3505
box -2 -3 34 103
use OAI22X1  OAI22X1_44
timestamp 1719641852
transform -1 0 2860 0 -1 3505
box -2 -3 42 103
use NAND2X1  NAND2X1_346
timestamp 1719641852
transform -1 0 2884 0 -1 3505
box -2 -3 26 103
use BUFX4  BUFX4_110
timestamp 1719641852
transform 1 0 2884 0 -1 3505
box -2 -3 34 103
use FILL  FILL_34_5_0
timestamp 1719641852
transform -1 0 2924 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_5_1
timestamp 1719641852
transform -1 0 2932 0 -1 3505
box -2 -3 10 103
use NAND2X1  NAND2X1_347
timestamp 1719641852
transform -1 0 2956 0 -1 3505
box -2 -3 26 103
use NAND2X1  NAND2X1_108
timestamp 1719641852
transform -1 0 2980 0 -1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_198
timestamp 1719641852
transform -1 0 3012 0 -1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_106
timestamp 1719641852
transform -1 0 3036 0 -1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_191
timestamp 1719641852
transform -1 0 3068 0 -1 3505
box -2 -3 34 103
use INVX1  INVX1_86
timestamp 1719641852
transform -1 0 3084 0 -1 3505
box -2 -3 18 103
use INVX8  INVX8_13
timestamp 1719641852
transform -1 0 3124 0 -1 3505
box -2 -3 42 103
use OR2X2  OR2X2_7
timestamp 1719641852
transform -1 0 3156 0 -1 3505
box -2 -3 34 103
use NOR2X1  NOR2X1_177
timestamp 1719641852
transform 1 0 3156 0 -1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_274
timestamp 1719641852
transform 1 0 3180 0 -1 3505
box -2 -3 34 103
use NAND3X1  NAND3X1_174
timestamp 1719641852
transform 1 0 3212 0 -1 3505
box -2 -3 34 103
use NAND3X1  NAND3X1_175
timestamp 1719641852
transform -1 0 3276 0 -1 3505
box -2 -3 34 103
use OAI21X1  OAI21X1_279
timestamp 1719641852
transform -1 0 3308 0 -1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_142
timestamp 1719641852
transform 1 0 3308 0 -1 3505
box -2 -3 26 103
use NAND3X1  NAND3X1_181
timestamp 1719641852
transform -1 0 3364 0 -1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_143
timestamp 1719641852
transform -1 0 3388 0 -1 3505
box -2 -3 26 103
use NOR2X1  NOR2X1_178
timestamp 1719641852
transform -1 0 3412 0 -1 3505
box -2 -3 26 103
use FILL  FILL_34_6_0
timestamp 1719641852
transform 1 0 3412 0 -1 3505
box -2 -3 10 103
use FILL  FILL_34_6_1
timestamp 1719641852
transform 1 0 3420 0 -1 3505
box -2 -3 10 103
use OR2X2  OR2X2_11
timestamp 1719641852
transform 1 0 3428 0 -1 3505
box -2 -3 34 103
use INVX2  INVX2_51
timestamp 1719641852
transform 1 0 3460 0 -1 3505
box -2 -3 18 103
use NAND2X1  NAND2X1_140
timestamp 1719641852
transform 1 0 3476 0 -1 3505
box -2 -3 26 103
use NAND2X1  NAND2X1_138
timestamp 1719641852
transform -1 0 3524 0 -1 3505
box -2 -3 26 103
use NAND3X1  NAND3X1_178
timestamp 1719641852
transform -1 0 3556 0 -1 3505
box -2 -3 34 103
use NAND3X1  NAND3X1_176
timestamp 1719641852
transform -1 0 3588 0 -1 3505
box -2 -3 34 103
use NAND3X1  NAND3X1_179
timestamp 1719641852
transform -1 0 3620 0 -1 3505
box -2 -3 34 103
use INVX8  INVX8_9
timestamp 1719641852
transform 1 0 3620 0 -1 3505
box -2 -3 42 103
use OAI21X1  OAI21X1_258
timestamp 1719641852
transform 1 0 3660 0 -1 3505
box -2 -3 34 103
use NAND3X1  NAND3X1_183
timestamp 1719641852
transform 1 0 3692 0 -1 3505
box -2 -3 34 103
use AOI21X1  AOI21X1_40
timestamp 1719641852
transform -1 0 3756 0 -1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_114
timestamp 1719641852
transform 1 0 3756 0 -1 3505
box -2 -3 26 103
use CLKBUF1  CLKBUF1_53
timestamp 1719641852
transform 1 0 4 0 1 3505
box -2 -3 74 103
use CLKBUF1  CLKBUF1_36
timestamp 1719641852
transform 1 0 76 0 1 3505
box -2 -3 74 103
use BUFX2  BUFX2_8
timestamp 1719641852
transform -1 0 172 0 1 3505
box -2 -3 26 103
use CLKBUF1  CLKBUF1_46
timestamp 1719641852
transform 1 0 172 0 1 3505
box -2 -3 74 103
use BUFX2  BUFX2_9
timestamp 1719641852
transform 1 0 244 0 1 3505
box -2 -3 26 103
use BUFX2  BUFX2_7
timestamp 1719641852
transform -1 0 292 0 1 3505
box -2 -3 26 103
use BUFX2  BUFX2_5
timestamp 1719641852
transform -1 0 316 0 1 3505
box -2 -3 26 103
use BUFX2  BUFX2_38
timestamp 1719641852
transform -1 0 340 0 1 3505
box -2 -3 26 103
use FILL  FILL_35_0_0
timestamp 1719641852
transform -1 0 348 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_0_1
timestamp 1719641852
transform -1 0 356 0 1 3505
box -2 -3 10 103
use DFFSR  DFFSR_67
timestamp 1719641852
transform -1 0 532 0 1 3505
box -2 -3 178 103
use BUFX2  BUFX2_42
timestamp 1719641852
transform -1 0 556 0 1 3505
box -2 -3 26 103
use DFFSR  DFFSR_71
timestamp 1719641852
transform -1 0 732 0 1 3505
box -2 -3 178 103
use BUFX2  BUFX2_4
timestamp 1719641852
transform 1 0 732 0 1 3505
box -2 -3 26 103
use BUFX2  BUFX2_53
timestamp 1719641852
transform -1 0 780 0 1 3505
box -2 -3 26 103
use FILL  FILL_35_1_0
timestamp 1719641852
transform -1 0 788 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_1_1
timestamp 1719641852
transform -1 0 796 0 1 3505
box -2 -3 10 103
use DFFSR  DFFSR_82
timestamp 1719641852
transform -1 0 972 0 1 3505
box -2 -3 178 103
use BUFX2  BUFX2_52
timestamp 1719641852
transform 1 0 972 0 1 3505
box -2 -3 26 103
use DFFSR  DFFSR_70
timestamp 1719641852
transform 1 0 996 0 1 3505
box -2 -3 178 103
use BUFX2  BUFX2_1
timestamp 1719641852
transform 1 0 1172 0 1 3505
box -2 -3 26 103
use BUFX2  BUFX2_41
timestamp 1719641852
transform 1 0 1196 0 1 3505
box -2 -3 26 103
use DFFSR  DFFSR_65
timestamp 1719641852
transform 1 0 1220 0 1 3505
box -2 -3 178 103
use FILL  FILL_35_2_0
timestamp 1719641852
transform 1 0 1396 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_2_1
timestamp 1719641852
transform 1 0 1404 0 1 3505
box -2 -3 10 103
use BUFX2  BUFX2_22
timestamp 1719641852
transform 1 0 1412 0 1 3505
box -2 -3 26 103
use BUFX2  BUFX2_24
timestamp 1719641852
transform 1 0 1436 0 1 3505
box -2 -3 26 103
use BUFX2  BUFX2_36
timestamp 1719641852
transform 1 0 1460 0 1 3505
box -2 -3 26 103
use BUFX2  BUFX2_23
timestamp 1719641852
transform 1 0 1484 0 1 3505
box -2 -3 26 103
use DFFSR  DFFSR_85
timestamp 1719641852
transform 1 0 1508 0 1 3505
box -2 -3 178 103
use BUFX2  BUFX2_56
timestamp 1719641852
transform 1 0 1684 0 1 3505
box -2 -3 26 103
use BUFX2  BUFX2_57
timestamp 1719641852
transform 1 0 1708 0 1 3505
box -2 -3 26 103
use DFFSR  DFFSR_88
timestamp 1719641852
transform 1 0 1732 0 1 3505
box -2 -3 178 103
use FILL  FILL_35_3_0
timestamp 1719641852
transform 1 0 1908 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_3_1
timestamp 1719641852
transform 1 0 1916 0 1 3505
box -2 -3 10 103
use BUFX2  BUFX2_59
timestamp 1719641852
transform 1 0 1924 0 1 3505
box -2 -3 26 103
use BUFX2  BUFX2_54
timestamp 1719641852
transform -1 0 1972 0 1 3505
box -2 -3 26 103
use AOI21X1  AOI21X1_269
timestamp 1719641852
transform -1 0 2004 0 1 3505
box -2 -3 34 103
use INVX4  INVX4_5
timestamp 1719641852
transform -1 0 2028 0 1 3505
box -2 -3 26 103
use CLKBUF1  CLKBUF1_27
timestamp 1719641852
transform -1 0 2100 0 1 3505
box -2 -3 74 103
use CLKBUF1  CLKBUF1_54
timestamp 1719641852
transform -1 0 2172 0 1 3505
box -2 -3 74 103
use NOR2X1  NOR2X1_346
timestamp 1719641852
transform 1 0 2172 0 1 3505
box -2 -3 26 103
use DFFSR  DFFSR_253
timestamp 1719641852
transform 1 0 2196 0 1 3505
box -2 -3 178 103
use NAND2X1  NAND2X1_345
timestamp 1719641852
transform -1 0 2396 0 1 3505
box -2 -3 26 103
use FILL  FILL_35_4_0
timestamp 1719641852
transform 1 0 2396 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_4_1
timestamp 1719641852
transform 1 0 2404 0 1 3505
box -2 -3 10 103
use NOR2X1  NOR2X1_349
timestamp 1719641852
transform 1 0 2412 0 1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_799
timestamp 1719641852
transform 1 0 2436 0 1 3505
box -2 -3 34 103
use AOI22X1  AOI22X1_85
timestamp 1719641852
transform -1 0 2508 0 1 3505
box -2 -3 42 103
use DFFSR  DFFSR_252
timestamp 1719641852
transform 1 0 2508 0 1 3505
box -2 -3 178 103
use DFFSR  DFFSR_250
timestamp 1719641852
transform 1 0 2684 0 1 3505
box -2 -3 178 103
use NOR2X1  NOR2X1_347
timestamp 1719641852
transform 1 0 2860 0 1 3505
box -2 -3 26 103
use NAND2X1  NAND2X1_344
timestamp 1719641852
transform 1 0 2884 0 1 3505
box -2 -3 26 103
use FILL  FILL_35_5_0
timestamp 1719641852
transform -1 0 2916 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_5_1
timestamp 1719641852
transform -1 0 2924 0 1 3505
box -2 -3 10 103
use OAI21X1  OAI21X1_796
timestamp 1719641852
transform -1 0 2956 0 1 3505
box -2 -3 34 103
use DFFSR  DFFSR_249
timestamp 1719641852
transform 1 0 2956 0 1 3505
box -2 -3 178 103
use NOR2X1  NOR2X1_48
timestamp 1719641852
transform 1 0 3132 0 1 3505
box -2 -3 26 103
use NAND2X1  NAND2X1_102
timestamp 1719641852
transform -1 0 3180 0 1 3505
box -2 -3 26 103
use OAI21X1  OAI21X1_795
timestamp 1719641852
transform -1 0 3212 0 1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_343
timestamp 1719641852
transform -1 0 3236 0 1 3505
box -2 -3 26 103
use INVX2  INVX2_42
timestamp 1719641852
transform -1 0 3252 0 1 3505
box -2 -3 18 103
use OAI21X1  OAI21X1_195
timestamp 1719641852
transform 1 0 3252 0 1 3505
box -2 -3 34 103
use AOI21X1  AOI21X1_46
timestamp 1719641852
transform 1 0 3284 0 1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_107
timestamp 1719641852
transform 1 0 3316 0 1 3505
box -2 -3 26 103
use AND2X2  AND2X2_18
timestamp 1719641852
transform -1 0 3372 0 1 3505
box -2 -3 34 103
use NAND2X1  NAND2X1_139
timestamp 1719641852
transform 1 0 3372 0 1 3505
box -2 -3 26 103
use NOR2X1  NOR2X1_176
timestamp 1719641852
transform -1 0 3420 0 1 3505
box -2 -3 26 103
use FILL  FILL_35_6_0
timestamp 1719641852
transform -1 0 3428 0 1 3505
box -2 -3 10 103
use FILL  FILL_35_6_1
timestamp 1719641852
transform -1 0 3436 0 1 3505
box -2 -3 10 103
use AOI21X1  AOI21X1_36
timestamp 1719641852
transform -1 0 3468 0 1 3505
box -2 -3 34 103
use NAND3X1  NAND3X1_180
timestamp 1719641852
transform 1 0 3468 0 1 3505
box -2 -3 34 103
use NOR2X1  NOR2X1_61
timestamp 1719641852
transform -1 0 3524 0 1 3505
box -2 -3 26 103
use INVX2  INVX2_49
timestamp 1719641852
transform 1 0 3524 0 1 3505
box -2 -3 18 103
use AND2X2  AND2X2_19
timestamp 1719641852
transform 1 0 3540 0 1 3505
box -2 -3 34 103
use NOR2X1  NOR2X1_60
timestamp 1719641852
transform -1 0 3596 0 1 3505
box -2 -3 26 103
use NOR2X1  NOR2X1_163
timestamp 1719641852
transform 1 0 3596 0 1 3505
box -2 -3 26 103
use BUFX4  BUFX4_197
timestamp 1719641852
transform -1 0 3652 0 1 3505
box -2 -3 34 103
use NAND3X1  NAND3X1_160
timestamp 1719641852
transform 1 0 3652 0 1 3505
box -2 -3 34 103
use BUFX4  BUFX4_194
timestamp 1719641852
transform -1 0 3716 0 1 3505
box -2 -3 34 103
use AND2X2  AND2X2_12
timestamp 1719641852
transform -1 0 3748 0 1 3505
box -2 -3 34 103
use FILL  FILL_36_1
timestamp 1719641852
transform 1 0 3748 0 1 3505
box -2 -3 10 103
use FILL  FILL_36_2
timestamp 1719641852
transform 1 0 3756 0 1 3505
box -2 -3 10 103
use FILL  FILL_36_3
timestamp 1719641852
transform 1 0 3764 0 1 3505
box -2 -3 10 103
use FILL  FILL_36_4
timestamp 1719641852
transform 1 0 3772 0 1 3505
box -2 -3 10 103
<< labels >>
flabel metal6 s 344 -30 360 -22 7 FreeSans 24 270 0 0 vdd
port 0 nsew
flabel metal6 s 848 -30 864 -22 7 FreeSans 24 270 0 0 gnd
port 1 nsew
flabel metal3 s -26 3138 -22 3142 7 FreeSans 24 0 0 0 wb_clk_i
port 2 nsew
flabel metal3 s -26 1338 -22 1342 7 FreeSans 24 0 0 0 wb_rst_i
port 3 nsew
flabel metal3 s -26 2538 -22 2542 7 FreeSans 24 0 0 0 wb_adr_i[0]
port 4 nsew
flabel metal2 s 2118 3628 2122 3632 3 FreeSans 24 90 0 0 wb_adr_i[1]
port 5 nsew
flabel metal3 s -26 1948 -22 1952 7 FreeSans 24 0 0 0 wb_adr_i[2]
port 6 nsew
flabel metal2 s 1462 3628 1466 3632 3 FreeSans 24 90 0 0 wb_adr_i[3]
port 7 nsew
flabel metal2 s 1382 3628 1386 3632 3 FreeSans 24 90 0 0 wb_adr_i[4]
port 8 nsew
flabel metal2 s 2062 3628 2066 3632 3 FreeSans 24 90 0 0 wb_dat_i[0]
port 9 nsew
flabel metal2 s 2230 3628 2234 3632 3 FreeSans 24 90 0 0 wb_dat_i[1]
port 10 nsew
flabel metal2 s 886 3628 890 3632 3 FreeSans 24 90 0 0 wb_dat_i[2]
port 11 nsew
flabel metal2 s 1270 3628 1274 3632 3 FreeSans 24 90 0 0 wb_dat_i[3]
port 12 nsew
flabel metal2 s 1334 3628 1338 3632 3 FreeSans 24 90 0 0 wb_dat_i[4]
port 13 nsew
flabel metal2 s 1974 3628 1978 3632 3 FreeSans 24 90 0 0 wb_dat_i[5]
port 14 nsew
flabel metal3 s -26 2648 -22 2652 7 FreeSans 24 0 0 0 wb_dat_i[6]
port 15 nsew
flabel metal3 s -26 2398 -22 2402 7 FreeSans 24 0 0 0 wb_dat_i[7]
port 16 nsew
flabel metal3 s -26 1848 -22 1852 7 FreeSans 24 0 0 0 wb_dat_i[8]
port 17 nsew
flabel metal3 s -26 1448 -22 1452 7 FreeSans 24 0 0 0 wb_dat_i[9]
port 18 nsew
flabel metal3 s -26 1168 -22 1172 7 FreeSans 24 0 0 0 wb_dat_i[10]
port 19 nsew
flabel metal2 s 1102 -22 1106 -18 7 FreeSans 24 270 0 0 wb_dat_i[11]
port 20 nsew
flabel metal3 s -26 1668 -22 1672 7 FreeSans 24 0 0 0 wb_dat_i[12]
port 21 nsew
flabel metal3 s -26 1648 -22 1652 7 FreeSans 24 0 0 0 wb_dat_i[13]
port 22 nsew
flabel metal3 s -26 1358 -22 1362 7 FreeSans 24 0 0 0 wb_dat_i[14]
port 23 nsew
flabel metal3 s -26 1148 -22 1152 7 FreeSans 24 0 0 0 wb_dat_i[15]
port 24 nsew
flabel metal2 s 2406 3628 2410 3632 3 FreeSans 24 90 0 0 wb_dat_i[16]
port 25 nsew
flabel metal2 s 2078 3628 2082 3632 3 FreeSans 24 90 0 0 wb_dat_i[17]
port 26 nsew
flabel metal2 s 1662 3628 1666 3632 3 FreeSans 24 90 0 0 wb_dat_i[18]
port 27 nsew
flabel metal2 s 1510 3628 1514 3632 3 FreeSans 24 90 0 0 wb_dat_i[19]
port 28 nsew
flabel metal2 s 1790 3628 1794 3632 3 FreeSans 24 90 0 0 wb_dat_i[20]
port 29 nsew
flabel metal2 s 1902 3628 1906 3632 3 FreeSans 24 90 0 0 wb_dat_i[21]
port 30 nsew
flabel metal2 s 1758 3628 1762 3632 3 FreeSans 24 90 0 0 wb_dat_i[22]
port 31 nsew
flabel metal2 s 1606 3628 1610 3632 3 FreeSans 24 90 0 0 wb_dat_i[23]
port 32 nsew
flabel metal2 s 1998 -22 2002 -18 7 FreeSans 24 270 0 0 wb_dat_i[24]
port 33 nsew
flabel metal2 s 1862 -22 1866 -18 7 FreeSans 24 270 0 0 wb_dat_i[25]
port 34 nsew
flabel metal2 s 1278 -22 1282 -18 7 FreeSans 24 270 0 0 wb_dat_i[26]
port 35 nsew
flabel metal2 s 2494 -22 2498 -18 7 FreeSans 24 270 0 0 wb_dat_i[27]
port 36 nsew
flabel metal2 s 2094 -22 2098 -18 7 FreeSans 24 270 0 0 wb_dat_i[28]
port 37 nsew
flabel metal2 s 1214 -22 1218 -18 7 FreeSans 24 270 0 0 wb_dat_i[29]
port 38 nsew
flabel metal2 s 1926 -22 1930 -18 7 FreeSans 24 270 0 0 wb_dat_i[30]
port 39 nsew
flabel metal2 s 1430 -22 1434 -18 7 FreeSans 24 270 0 0 wb_dat_i[31]
port 40 nsew
flabel metal2 s 958 3628 962 3632 3 FreeSans 24 90 0 0 wb_sel_i[0]
port 41 nsew
flabel metal3 s -26 1548 -22 1552 7 FreeSans 24 0 0 0 wb_sel_i[1]
port 42 nsew
flabel metal2 s 1774 3628 1778 3632 3 FreeSans 24 90 0 0 wb_sel_i[2]
port 43 nsew
flabel metal2 s 1238 -22 1242 -18 7 FreeSans 24 270 0 0 wb_sel_i[3]
port 44 nsew
flabel metal2 s 270 -22 274 -18 7 FreeSans 24 270 0 0 wb_we_i
port 45 nsew
flabel metal2 s 254 -22 258 -18 7 FreeSans 24 270 0 0 wb_stb_i
port 46 nsew
flabel metal2 s 238 -22 242 -18 7 FreeSans 24 270 0 0 wb_cyc_i
port 47 nsew
flabel metal3 s 3806 1448 3810 1452 3 FreeSans 24 0 0 0 miso_pad_i
port 48 nsew
flabel metal2 s 1478 3628 1482 3632 3 FreeSans 24 90 0 0 wb_dat_o[0]
port 49 nsew
flabel metal3 s -26 3248 -22 3252 7 FreeSans 24 0 0 0 wb_dat_o[1]
port 50 nsew
flabel metal2 s 326 3628 330 3632 3 FreeSans 24 90 0 0 wb_dat_o[2]
port 51 nsew
flabel metal2 s 1070 3628 1074 3632 3 FreeSans 24 90 0 0 wb_dat_o[3]
port 52 nsew
flabel metal3 s -26 2558 -22 2562 7 FreeSans 24 0 0 0 wb_dat_o[4]
port 53 nsew
flabel metal2 s 1206 3628 1210 3632 3 FreeSans 24 90 0 0 wb_dat_o[5]
port 54 nsew
flabel metal2 s 542 3628 546 3632 3 FreeSans 24 90 0 0 wb_dat_o[6]
port 55 nsew
flabel metal3 s -26 2368 -22 2372 7 FreeSans 24 0 0 0 wb_dat_o[7]
port 56 nsew
flabel metal3 s -26 1968 -22 1972 7 FreeSans 24 0 0 0 wb_dat_o[8]
port 57 nsew
flabel metal3 s -26 2348 -22 2352 7 FreeSans 24 0 0 0 wb_dat_o[9]
port 58 nsew
flabel metal3 s -26 1378 -22 1382 7 FreeSans 24 0 0 0 wb_dat_o[10]
port 59 nsew
flabel metal3 s -26 1748 -22 1752 7 FreeSans 24 0 0 0 wb_dat_o[11]
port 60 nsew
flabel metal2 s 214 3628 218 3632 3 FreeSans 24 90 0 0 wb_dat_o[12]
port 61 nsew
flabel metal3 s -26 1588 -22 1592 7 FreeSans 24 0 0 0 wb_dat_o[13]
port 62 nsew
flabel metal2 s 1254 -22 1258 -18 7 FreeSans 24 270 0 0 wb_dat_o[14]
port 63 nsew
flabel metal2 s 630 -22 634 -18 7 FreeSans 24 270 0 0 wb_dat_o[15]
port 64 nsew
flabel metal2 s 982 3628 986 3632 3 FreeSans 24 90 0 0 wb_dat_o[16]
port 65 nsew
flabel metal2 s 766 3628 770 3632 3 FreeSans 24 90 0 0 wb_dat_o[17]
port 66 nsew
flabel metal2 s 1958 3628 1962 3632 3 FreeSans 24 90 0 0 wb_dat_o[18]
port 67 nsew
flabel metal3 s -26 2468 -22 2472 7 FreeSans 24 0 0 0 wb_dat_o[19]
port 68 nsew
flabel metal2 s 1694 3628 1698 3632 3 FreeSans 24 90 0 0 wb_dat_o[20]
port 69 nsew
flabel metal2 s 1718 3628 1722 3632 3 FreeSans 24 90 0 0 wb_dat_o[21]
port 70 nsew
flabel metal3 s -26 2748 -22 2752 7 FreeSans 24 0 0 0 wb_dat_o[22]
port 71 nsew
flabel metal2 s 1934 3628 1938 3632 3 FreeSans 24 90 0 0 wb_dat_o[23]
port 72 nsew
flabel metal2 s 1022 -22 1026 -18 7 FreeSans 24 270 0 0 wb_dat_o[24]
port 73 nsew
flabel metal2 s 1534 -22 1538 -18 7 FreeSans 24 270 0 0 wb_dat_o[25]
port 74 nsew
flabel metal3 s -26 48 -22 52 7 FreeSans 24 270 0 0 wb_dat_o[26]
port 75 nsew
flabel metal2 s 1734 -22 1738 -18 7 FreeSans 24 270 0 0 wb_dat_o[27]
port 76 nsew
flabel metal2 s 182 -22 186 -18 7 FreeSans 24 270 0 0 wb_dat_o[28]
port 77 nsew
flabel metal2 s 1446 -22 1450 -18 7 FreeSans 24 270 0 0 wb_dat_o[29]
port 78 nsew
flabel metal2 s 382 -22 386 -18 7 FreeSans 24 270 0 0 wb_dat_o[30]
port 79 nsew
flabel metal2 s 214 -22 218 -18 7 FreeSans 24 270 0 0 wb_dat_o[31]
port 80 nsew
flabel metal3 s -26 3368 -22 3372 7 FreeSans 24 0 0 0 wb_ack_o
port 81 nsew
flabel metal3 s -26 148 -22 152 7 FreeSans 24 0 0 0 wb_err_o
port 82 nsew
flabel metal3 s -26 3348 -22 3352 7 FreeSans 24 0 0 0 wb_int_o
port 83 nsew
flabel metal2 s 430 3628 434 3632 3 FreeSans 24 90 0 0 ss_pad_o[0]
port 84 nsew
flabel metal2 s 742 3628 746 3632 3 FreeSans 24 90 0 0 ss_pad_o[1]
port 85 nsew
flabel metal2 s 302 3628 306 3632 3 FreeSans 24 90 0 0 ss_pad_o[2]
port 86 nsew
flabel metal3 s -26 2868 -22 2872 7 FreeSans 24 0 0 0 ss_pad_o[3]
port 87 nsew
flabel metal2 s 278 3628 282 3632 3 FreeSans 24 90 0 0 ss_pad_o[4]
port 88 nsew
flabel metal2 s 158 3628 162 3632 3 FreeSans 24 90 0 0 ss_pad_o[5]
port 89 nsew
flabel metal2 s 254 3628 258 3632 3 FreeSans 24 90 0 0 ss_pad_o[6]
port 90 nsew
flabel metal3 s -26 2448 -22 2452 7 FreeSans 24 0 0 0 ss_pad_o[7]
port 91 nsew
flabel metal3 s -26 2248 -22 2252 7 FreeSans 24 0 0 0 ss_pad_o[8]
port 92 nsew
flabel metal3 s -26 2148 -22 2152 7 FreeSans 24 0 0 0 ss_pad_o[9]
port 93 nsew
flabel metal3 s -26 1068 -22 1072 7 FreeSans 24 0 0 0 ss_pad_o[10]
port 94 nsew
flabel metal3 s -26 1988 -22 1992 7 FreeSans 24 0 0 0 ss_pad_o[11]
port 95 nsew
flabel metal3 s -26 2048 -22 2052 7 FreeSans 24 0 0 0 ss_pad_o[12]
port 96 nsew
flabel metal3 s -26 2068 -22 2072 7 FreeSans 24 0 0 0 ss_pad_o[13]
port 97 nsew
flabel metal3 s -26 2848 -22 2852 7 FreeSans 24 0 0 0 ss_pad_o[14]
port 98 nsew
flabel metal3 s -26 1048 -22 1052 7 FreeSans 24 0 0 0 ss_pad_o[15]
port 99 nsew
flabel metal2 s 1174 3628 1178 3632 3 FreeSans 24 90 0 0 ss_pad_o[16]
port 100 nsew
flabel metal3 s -26 3048 -22 3052 7 FreeSans 24 0 0 0 ss_pad_o[17]
port 101 nsew
flabel metal2 s 1574 3628 1578 3632 3 FreeSans 24 90 0 0 ss_pad_o[18]
port 102 nsew
flabel metal2 s 1422 3628 1426 3632 3 FreeSans 24 90 0 0 ss_pad_o[19]
port 103 nsew
flabel metal2 s 1526 3628 1530 3632 3 FreeSans 24 90 0 0 ss_pad_o[20]
port 104 nsew
flabel metal2 s 1446 3628 1450 3632 3 FreeSans 24 90 0 0 ss_pad_o[21]
port 105 nsew
flabel metal3 s -26 2948 -22 2952 7 FreeSans 24 0 0 0 ss_pad_o[22]
port 106 nsew
flabel metal3 s -26 3448 -22 3452 7 FreeSans 24 0 0 0 ss_pad_o[23]
port 107 nsew
flabel metal2 s 582 -22 586 -18 7 FreeSans 24 270 0 0 ss_pad_o[24]
port 108 nsew
flabel metal2 s 766 -22 770 -18 7 FreeSans 24 270 0 0 ss_pad_o[25]
port 109 nsew
flabel metal2 s 294 -22 298 -18 7 FreeSans 24 270 0 0 ss_pad_o[26]
port 110 nsew
flabel metal2 s 366 -22 370 -18 7 FreeSans 24 270 0 0 ss_pad_o[27]
port 111 nsew
flabel metal2 s 726 -22 730 -18 7 FreeSans 24 270 0 0 ss_pad_o[28]
port 112 nsew
flabel metal2 s 606 -22 610 -18 7 FreeSans 24 270 0 0 ss_pad_o[29]
port 113 nsew
flabel metal2 s 678 -22 682 -18 7 FreeSans 24 270 0 0 ss_pad_o[30]
port 114 nsew
flabel metal2 s 318 -22 322 -18 7 FreeSans 24 270 0 0 ss_pad_o[31]
port 115 nsew
flabel metal3 s -26 1568 -22 1572 7 FreeSans 24 0 0 0 sclk_pad_o
port 116 nsew
flabel metal2 s 1190 3628 1194 3632 3 FreeSans 24 90 0 0 mosi_pad_o
port 117 nsew
<< end >>
