* NGSPICE file created from spi_top.ext - technology: scmos

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for DFFSR abstract view
.subckt DFFSR Q CLK R S D gnd vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for OAI22X1 abstract view
.subckt OAI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX4 abstract view
.subckt BUFX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for XNOR2X1 abstract view
.subckt XNOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX8 abstract view
.subckt INVX8 A gnd Y vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for NOR3X1 abstract view
.subckt NOR3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 A gnd Y vdd
.ends

* Black-box entry subcircuit for MUX2X1 abstract view
.subckt MUX2X1 A B S gnd Y vdd
.ends

* Black-box entry subcircuit for XOR2X1 abstract view
.subckt XOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX4 abstract view
.subckt INVX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

.subckt spi_top vdd gnd wb_clk_i wb_rst_i wb_adr_i[0] wb_adr_i[1] wb_adr_i[2] wb_adr_i[3]
+ wb_adr_i[4] wb_dat_i[0] wb_dat_i[1] wb_dat_i[2] wb_dat_i[3] wb_dat_i[4] wb_dat_i[5]
+ wb_dat_i[6] wb_dat_i[7] wb_dat_i[8] wb_dat_i[9] wb_dat_i[10] wb_dat_i[11] wb_dat_i[12]
+ wb_dat_i[13] wb_dat_i[14] wb_dat_i[15] wb_dat_i[16] wb_dat_i[17] wb_dat_i[18] wb_dat_i[19]
+ wb_dat_i[20] wb_dat_i[21] wb_dat_i[22] wb_dat_i[23] wb_dat_i[24] wb_dat_i[25] wb_dat_i[26]
+ wb_dat_i[27] wb_dat_i[28] wb_dat_i[29] wb_dat_i[30] wb_dat_i[31] wb_sel_i[0] wb_sel_i[1]
+ wb_sel_i[2] wb_sel_i[3] wb_we_i wb_stb_i wb_cyc_i miso_pad_i wb_dat_o[0] wb_dat_o[1]
+ wb_dat_o[2] wb_dat_o[3] wb_dat_o[4] wb_dat_o[5] wb_dat_o[6] wb_dat_o[7] wb_dat_o[8]
+ wb_dat_o[9] wb_dat_o[10] wb_dat_o[11] wb_dat_o[12] wb_dat_o[13] wb_dat_o[14] wb_dat_o[15]
+ wb_dat_o[16] wb_dat_o[17] wb_dat_o[18] wb_dat_o[19] wb_dat_o[20] wb_dat_o[21] wb_dat_o[22]
+ wb_dat_o[23] wb_dat_o[24] wb_dat_o[25] wb_dat_o[26] wb_dat_o[27] wb_dat_o[28] wb_dat_o[29]
+ wb_dat_o[30] wb_dat_o[31] wb_ack_o wb_err_o wb_int_o ss_pad_o[0] ss_pad_o[1] ss_pad_o[2]
+ ss_pad_o[3] ss_pad_o[4] ss_pad_o[5] ss_pad_o[6] ss_pad_o[7] ss_pad_o[8] ss_pad_o[9]
+ ss_pad_o[10] ss_pad_o[11] ss_pad_o[12] ss_pad_o[13] ss_pad_o[14] ss_pad_o[15] ss_pad_o[16]
+ ss_pad_o[17] ss_pad_o[18] ss_pad_o[19] ss_pad_o[20] ss_pad_o[21] ss_pad_o[22] ss_pad_o[23]
+ ss_pad_o[24] ss_pad_o[25] ss_pad_o[26] ss_pad_o[27] ss_pad_o[28] ss_pad_o[29] ss_pad_o[30]
+ ss_pad_o[31] sclk_pad_o mosi_pad_o
XFILL_9_6_0 gnd vdd FILL
XFILL_17_5_0 gnd vdd FILL
XOAI21X1_360 OAI21X1_360/A OAI21X1_359/Y OAI21X1_356/Y gnd DFFSR_234/D vdd OAI21X1
XOAI21X1_371 NOR2X1_215/Y INVX2_77/Y BUFX4_51/Y gnd AOI21X1_119/C vdd OAI21X1
XAND2X2_5 AND2X2_5/A AND2X2_5/B gnd AND2X2_5/Y vdd AND2X2
XOAI21X1_382 BUFX4_67/Y NAND2X1_230/Y AOI21X1_124/Y gnd AOI21X1_126/B vdd OAI21X1
XOAI21X1_393 OAI21X1_393/A OAI21X1_392/Y OAI21X1_389/Y gnd DFFSR_224/D vdd OAI21X1
XFILL_32_3_0 gnd vdd FILL
XFILL_23_3_0 gnd vdd FILL
XFILL_6_4_0 gnd vdd FILL
XFILL_14_3_0 gnd vdd FILL
XOAI21X1_190 INVX2_18/A NAND2X1_104/Y OAI21X1_190/C gnd INVX2_47/A vdd OAI21X1
XDFFSR_9 INVX2_1/A DFFSR_9/CLK DFFSR_9/R vdd DFFSR_9/D gnd vdd DFFSR
XNAND2X1_10 BUFX4_161/Y wb_dat_i[17] gnd OAI21X1_19/C vdd NAND2X1
XNAND2X1_43 AOI21X1_5/Y NOR2X1_8/Y gnd DFFSR_69/D vdd NAND2X1
XNAND2X1_32 BUFX4_85/Y wb_dat_i[7] gnd OAI21X1_92/C vdd NAND2X1
XNAND2X1_21 BUFX4_5/Y wb_dat_i[12] gnd OAI21X1_71/C vdd NAND2X1
XNAND2X1_65 DFFSR_137/Q AOI21X1_1/B gnd NAND3X1_91/B vdd NAND2X1
XNAND2X1_54 AOI21X1_12/Y NOR2X1_15/Y gnd DFFSR_76/D vdd NAND2X1
XNAND2X1_87 OR2X2_2/B BUFX4_1/Y gnd NAND2X1_87/Y vdd NAND2X1
XNAND2X1_76 wb_stb_i wb_cyc_i gnd NOR2X1_18/B vdd NAND2X1
XNAND2X1_98 AND2X2_8/B AND2X2_8/A gnd OR2X2_5/A vdd NAND2X1
XAOI21X1_269 AOI22X1_85/D AOI22X1_85/C NOR2X1_350/Y gnd DFFSR_245/D vdd AOI21X1
XAOI21X1_203 AOI21X1_202/Y AOI21X1_203/B NOR2X1_275/Y gnd DFFSR_169/D vdd AOI21X1
XAOI21X1_236 AOI21X1_235/Y OAI21X1_636/Y NOR2X1_291/Y gnd DFFSR_152/D vdd AOI21X1
XAOI22X1_41 AOI22X1_41/A NOR2X1_189/Y INVX2_164/A AOI22X1_41/D gnd AOI21X1_67/A vdd
+ AOI22X1
XAOI22X1_30 BUFX4_21/Y INVX1_7/A INVX2_65/A INVX8_6/Y gnd AOI22X1_30/Y vdd AOI22X1
XAOI21X1_247 INVX1_97/A INVX1_156/Y BUFX4_212/Y gnd AOI22X1_82/D vdd AOI21X1
XAOI21X1_225 AOI21X1_225/A OAI21X1_622/Y NOR2X1_286/Y gnd DFFSR_158/D vdd AOI21X1
XAOI21X1_258 INVX2_123/Y AOI21X1_258/B BUFX4_34/Y gnd OAI21X1_769/C vdd AOI21X1
XAOI21X1_214 BUFX4_34/Y AOI21X1_214/B BUFX4_210/Y gnd AOI21X1_215/A vdd AOI21X1
XAOI22X1_85 AOI22X1_85/A AND2X2_33/Y AOI22X1_85/C AOI22X1_85/D gnd AOI22X1_85/Y vdd
+ AOI22X1
XAOI22X1_52 AOI22X1_52/A AOI21X1_79/Y AOI21X1_80/Y AOI22X1_52/D gnd AOI22X1_52/Y vdd
+ AOI22X1
XAOI22X1_74 INVX2_68/A INVX4_9/A INVX4_8/A INVX2_72/A gnd AOI22X1_74/Y vdd AOI22X1
XAOI22X1_63 DFFSR_239/Q INVX8_14/A INVX4_8/A INVX1_53/A gnd AOI22X1_63/Y vdd AOI22X1
XNAND3X1_207 OAI21X1_310/Y NAND3X1_207/B AOI22X1_66/Y gnd AOI22X1_68/A vdd NAND3X1
XOAI22X1_3 BUFX4_78/Y INVX2_10/Y INVX1_28/Y OAI22X1_1/D gnd NOR2X1_5/A vdd OAI22X1
XFILL_30_6_1 gnd vdd FILL
XDFFSR_216 INVX1_37/A DFFSR_36/CLK DFFSR_198/R vdd DFFSR_216/D gnd vdd DFFSR
XDFFSR_205 DFFSR_205/Q CLKBUF1_33/Y DFFSR_194/R vdd DFFSR_205/D gnd vdd DFFSR
XDFFSR_249 INVX2_48/A CLKBUF1_37/Y DFFSR_165/R vdd DFFSR_249/D gnd vdd DFFSR
XDFFSR_238 INVX2_67/A CLKBUF1_24/Y DFFSR_194/R vdd DFFSR_238/D gnd vdd DFFSR
XDFFSR_227 INVX1_62/A DFFSR_92/CLK DFFSR_236/R vdd DFFSR_227/D gnd vdd DFFSR
XFILL_21_6_1 gnd vdd FILL
XFILL_20_1_0 gnd vdd FILL
XINVX2_45 INVX2_45/A gnd INVX2_45/Y vdd INVX2
XINVX2_78 INVX2_78/A gnd INVX2_78/Y vdd INVX2
XINVX2_56 INVX2_56/A gnd INVX2_56/Y vdd INVX2
XINVX2_12 DFFSR_4/Q gnd INVX2_12/Y vdd INVX2
XINVX2_34 OR2X2_2/A gnd INVX2_34/Y vdd INVX2
XINVX2_23 DFFSR_55/Q gnd INVX2_23/Y vdd INVX2
XINVX2_67 INVX2_67/A gnd INVX2_67/Y vdd INVX2
XFILL_28_2_0 gnd vdd FILL
XINVX2_89 INVX2_89/A gnd INVX2_89/Y vdd INVX2
XFILL_3_2_0 gnd vdd FILL
XOAI21X1_19 INVX1_10/Y BUFX4_162/Y OAI21X1_19/C gnd NAND3X1_12/B vdd OAI21X1
XFILL_11_1_0 gnd vdd FILL
XFILL_12_6_1 gnd vdd FILL
XFILL_19_2_0 gnd vdd FILL
XNAND2X1_239 wb_dat_i[6] BUFX4_79/Y gnd NAND2X1_239/Y vdd NAND2X1
XNAND2X1_228 INVX8_14/A INVX1_129/Y gnd AOI21X1_121/B vdd NAND2X1
XNAND2X1_217 INVX1_126/Y NOR2X1_190/Y gnd INVX1_127/A vdd NAND2X1
XNAND2X1_206 BUFX4_71/Y wb_dat_i[27] gnd OAI21X1_567/C vdd NAND2X1
XBUFX4_190 BUFX4_193/A gnd BUFX4_190/Y vdd BUFX4
XNOR2X1_294 OR2X2_17/B NOR2X1_310/B gnd NOR2X1_294/Y vdd NOR2X1
XNOR2X1_250 INVX4_7/Y INVX1_136/Y gnd NOR2X1_250/Y vdd NOR2X1
XOAI21X1_712 BUFX4_60/Y OAI21X1_712/B OAI21X1_711/Y gnd OAI21X1_714/A vdd OAI21X1
XNOR2X1_261 INVX4_8/Y OR2X2_15/A gnd NOR2X1_261/Y vdd NOR2X1
XOAI21X1_723 INVX1_151/A OR2X2_18/B INVX2_117/Y gnd OAI21X1_724/C vdd OAI21X1
XOAI21X1_701 BUFX4_64/Y OR2X2_18/Y OAI21X1_700/Y gnd OAI21X1_702/A vdd OAI21X1
XNOR2X1_272 INVX4_9/Y NOR2X1_287/B gnd NOR2X1_272/Y vdd NOR2X1
XNOR2X1_283 INVX2_61/A BUFX4_118/Y gnd NOR2X1_283/Y vdd NOR2X1
XOAI21X1_734 NOR2X1_324/Y OAI21X1_733/Y NAND2X1_326/Y gnd DFFSR_116/D vdd OAI21X1
XOAI21X1_767 AOI21X1_256/Y OAI21X1_766/Y OAI21X1_763/Y gnd DFFSR_187/D vdd OAI21X1
XOAI21X1_789 BUFX4_60/Y OAI21X1_789/B OAI21X1_788/Y gnd OAI21X1_790/A vdd OAI21X1
XOAI21X1_778 BUFX4_59/Y OR2X2_21/Y OAI21X1_778/C gnd AOI21X1_267/B vdd OAI21X1
XOAI21X1_745 AOI21X1_250/Y OAI21X1_744/Y OAI21X1_741/Y gnd DFFSR_227/D vdd OAI21X1
XOAI21X1_756 NOR2X1_329/Y INVX2_124/Y BUFX4_167/Y gnd AOI21X1_253/C vdd OAI21X1
XBUFX4_85 wb_sel_i[0] gnd BUFX4_85/Y vdd BUFX4
XBUFX4_52 BUFX4_52/A gnd BUFX4_52/Y vdd BUFX4
XBUFX4_74 wb_sel_i[3] gnd MUX2X1_6/S vdd BUFX4
XBUFX4_41 BUFX4_45/A gnd BUFX4_41/Y vdd BUFX4
XBUFX4_63 BUFX4_61/A gnd BUFX4_63/Y vdd BUFX4
XBUFX4_96 BUFX4_98/A gnd BUFX4_96/Y vdd BUFX4
XBUFX4_30 BUFX4_32/A gnd BUFX4_30/Y vdd BUFX4
XFILL_35_5_1 gnd vdd FILL
XFILL_34_0_0 gnd vdd FILL
XOR2X2_11 OR2X2_11/A INVX2_49/Y gnd OR2X2_11/Y vdd OR2X2
XOR2X2_4 OR2X2_4/A OR2X2_4/B gnd OR2X2_4/Y vdd OR2X2
XXNOR2X1_6 XOR2X1_2/A XOR2X1_2/B gnd XNOR2X1_6/Y vdd XNOR2X1
XFILL_26_5_1 gnd vdd FILL
XFILL_25_0_0 gnd vdd FILL
XFILL_1_5_1 gnd vdd FILL
XFILL_0_0_0 gnd vdd FILL
XOAI21X1_553 BUFX4_211/Y BUFX4_28/Y DFFSR_180/Q gnd OAI21X1_553/Y vdd OAI21X1
XOAI21X1_542 AOI21X1_185/Y OAI21X1_541/Y OAI21X1_542/C gnd DFFSR_183/D vdd OAI21X1
XOAI21X1_531 BUFX4_169/Y OAI21X1_531/B BUFX4_37/Y gnd OAI21X1_532/B vdd OAI21X1
XINVX8_22 INVX8_22/A gnd INVX8_22/Y vdd INVX8
XINVX1_6 INVX1_6/A gnd INVX1_6/Y vdd INVX1
XOAI21X1_564 BUFX4_63/Y NAND2X1_259/Y OAI21X1_564/C gnd AOI21X1_195/B vdd OAI21X1
XINVX8_11 INVX8_11/A gnd INVX8_11/Y vdd INVX8
XOAI21X1_520 INVX2_98/Y BUFX4_7/Y NAND2X1_238/Y gnd OAI21X1_521/B vdd OAI21X1
XOAI21X1_575 BUFX4_99/Y INVX8_11/Y AND2X2_24/A gnd NOR2X1_287/B vdd OAI21X1
XOAI21X1_586 NOR2X1_274/Y INVX2_54/Y BUFX4_121/Y gnd AOI21X1_200/C vdd OAI21X1
XOAI21X1_597 BUFX4_98/Y INVX8_11/Y INVX1_136/A gnd NOR2X1_280/B vdd OAI21X1
XFILL_9_6_1 gnd vdd FILL
XFILL_8_1_0 gnd vdd FILL
XFILL_17_5_1 gnd vdd FILL
XFILL_16_0_0 gnd vdd FILL
XOAI21X1_372 INVX2_77/Y BUFX4_163/Y NAND2X1_224/Y gnd OAI21X1_373/B vdd OAI21X1
XOAI21X1_361 BUFX4_221/Y INVX8_19/A DFFSR_233/Q gnd OAI21X1_365/C vdd OAI21X1
XOAI21X1_350 OAI21X1_350/A OAI21X1_349/Y OAI21X1_350/C gnd DFFSR_237/D vdd OAI21X1
XOAI21X1_394 BUFX4_67/Y NAND2X1_234/Y OAI21X1_394/C gnd AOI21X1_131/B vdd OAI21X1
XOAI21X1_383 INVX2_62/Y BUFX4_12/Y NAND2X1_231/Y gnd OAI21X1_383/Y vdd OAI21X1
XAND2X2_6 AND2X2_6/A AND2X2_6/B gnd AND2X2_6/Y vdd AND2X2
XFILL_32_3_1 gnd vdd FILL
XFILL_23_3_1 gnd vdd FILL
XFILL_6_4_1 gnd vdd FILL
XFILL_14_3_1 gnd vdd FILL
XOAI21X1_191 OR2X2_8/Y INVX2_43/A INVX2_48/A gnd NAND2X1_106/A vdd OAI21X1
XAOI22X1_1 DFFSR_164/Q AOI22X1_1/B INVX8_5/Y DFFSR_196/Q gnd AOI22X1_1/Y vdd AOI22X1
XOAI21X1_180 OAI21X1_179/Y INVX1_77/Y OAI21X1_180/C gnd DFFSR_115/D vdd OAI21X1
XNAND2X1_33 BUFX4_103/Y OR2X2_3/B gnd NAND2X1_33/Y vdd NAND2X1
XNAND2X1_77 INVX1_19/A INVX4_11/A gnd OAI22X1_39/D vdd NAND2X1
XNAND2X1_11 BUFX4_163/Y wb_dat_i[18] gnd OAI21X1_21/C vdd NAND2X1
XNAND2X1_66 INVX2_56/A AOI21X1_1/B gnd NAND3X1_92/A vdd NAND2X1
XNAND2X1_44 AOI21X1_6/Y NOR2X1_9/Y gnd DFFSR_70/D vdd NAND2X1
XNAND2X1_55 NAND3X1_84/Y NAND2X1_55/B gnd AOI21X1_13/C vdd NAND2X1
XNAND2X1_22 BUFX4_7/Y wb_dat_i[13] gnd OAI21X1_73/C vdd NAND2X1
XNAND2X1_88 INVX2_32/A BUFX4_1/Y gnd NAND2X1_88/Y vdd NAND2X1
XNAND2X1_99 INVX1_76/Y AND2X2_8/A gnd OR2X2_6/A vdd NAND2X1
XAOI22X1_42 AOI22X1_42/A AOI21X1_60/Y AOI22X1_42/C INVX1_117/Y gnd AOI22X1_42/Y vdd
+ AOI22X1
XAOI21X1_237 INVX2_115/Y AOI21X1_237/B BUFX4_33/Y gnd OAI21X1_638/C vdd AOI21X1
XAOI21X1_204 INVX2_88/Y NAND2X1_265/Y BUFX4_31/Y gnd OAI21X1_593/C vdd AOI21X1
XAOI22X1_20 BUFX4_21/Y INVX1_2/A INVX2_141/A INVX8_6/Y gnd NAND3X1_95/C vdd AOI22X1
XAOI22X1_31 INVX2_126/A BUFX4_127/Y INVX8_5/Y INVX2_127/A gnd AOI22X1_31/Y vdd AOI22X1
XAOI22X1_75 INVX1_51/A INVX4_10/A INVX8_22/A INVX1_93/A gnd AOI22X1_75/Y vdd AOI22X1
XAOI21X1_248 INVX1_94/A INVX1_157/Y BUFX4_210/Y gnd AOI22X1_83/D vdd AOI21X1
XAOI22X1_64 INVX1_52/A INVX4_10/A INVX8_22/A INVX1_96/A gnd AOI22X1_64/Y vdd AOI22X1
XAOI21X1_259 BUFX4_34/Y AOI21X1_259/B BUFX4_210/Y gnd AOI21X1_259/Y vdd AOI21X1
XAOI21X1_215 AOI21X1_215/A AOI21X1_215/B NOR2X1_283/Y gnd DFFSR_162/D vdd AOI21X1
XAOI22X1_53 AOI22X1_53/A AOI22X1_53/B AOI21X1_82/Y AOI22X1_53/D gnd AOI22X1_53/Y vdd
+ AOI22X1
XAOI21X1_226 NOR2X1_287/Y BUFX4_64/Y AOI21X1_226/C gnd OAI21X1_627/A vdd AOI21X1
XNAND3X1_208 NAND3X1_208/A OAI21X1_313/Y AOI22X1_67/Y gnd AOI22X1_68/D vdd NAND3X1
XOAI22X1_4 OAI22X1_4/A INVX2_32/Y OAI22X1_4/C INVX1_29/Y gnd NOR2X1_5/B vdd OAI22X1
XDFFSR_228 AOI22X1_2/C CLKBUF1_12/Y BUFX4_130/Y vdd DFFSR_228/D gnd vdd DFFSR
XDFFSR_239 DFFSR_239/Q CLKBUF1_32/A DFFSR_236/R vdd DFFSR_239/D gnd vdd DFFSR
XDFFSR_206 INVX2_69/A DFFSR_26/CLK DFFSR_174/R vdd DFFSR_206/D gnd vdd DFFSR
XDFFSR_217 INVX1_40/A CLKBUF1_45/Y DFFSR_167/R vdd DFFSR_217/D gnd vdd DFFSR
XFILL_20_1_1 gnd vdd FILL
XINVX2_46 INVX2_46/A gnd INVX2_46/Y vdd INVX2
XINVX2_13 DFFSR_5/Q gnd INVX2_13/Y vdd INVX2
XINVX2_35 DFFSR_51/Q gnd INVX2_35/Y vdd INVX2
XINVX2_79 INVX2_79/A gnd INVX2_79/Y vdd INVX2
XINVX2_57 INVX1_43/A gnd INVX2_57/Y vdd INVX2
XINVX2_68 INVX2_68/A gnd INVX2_68/Y vdd INVX2
XINVX2_24 INVX2_24/A gnd INVX2_24/Y vdd INVX2
XFILL_28_2_1 gnd vdd FILL
XFILL_3_2_1 gnd vdd FILL
XFILL_11_1_1 gnd vdd FILL
XFILL_19_2_1 gnd vdd FILL
XNAND2X1_229 NAND2X1_9/B wb_dat_i[16] gnd NAND2X1_229/Y vdd NAND2X1
XNAND2X1_218 INVX8_14/A INVX1_127/Y gnd NAND2X1_218/Y vdd NAND2X1
XNAND2X1_207 INVX1_122/A NOR2X1_191/Y gnd NOR2X1_238/B vdd NAND2X1
XBUFX4_191 BUFX4_193/A gnd AOI21X1_2/B vdd BUFX4
XNOR2X1_251 BUFX4_152/Y OR2X2_13/B gnd INVX1_137/A vdd NOR2X1
XNOR2X1_240 DFFSR_205/Q BUFX4_35/Y gnd NOR2X1_240/Y vdd NOR2X1
XBUFX4_180 AND2X2_1/Y gnd BUFX4_180/Y vdd BUFX4
XNOR2X1_295 OR2X2_17/B NOR2X1_282/B gnd NOR2X1_295/Y vdd NOR2X1
XOAI21X1_713 INVX2_60/Y BUFX4_83/Y NAND2X1_239/Y gnd NAND2X1_315/B vdd OAI21X1
XNOR2X1_262 INVX4_8/Y NOR2X1_262/B gnd NOR2X1_262/Y vdd NOR2X1
XOAI21X1_724 BUFX4_96/Y INVX1_132/Y OAI21X1_724/C gnd OAI21X1_725/B vdd OAI21X1
XOAI21X1_702 OAI21X1_702/A BUFX4_208/Y NAND2X1_308/Y gnd DFFSR_128/D vdd OAI21X1
XOAI21X1_735 BUFX4_205/Y BUFX4_29/Y INVX2_127/A gnd OAI21X1_735/Y vdd OAI21X1
XOAI21X1_757 INVX2_124/Y BUFX4_8/Y NAND2X1_328/Y gnd OAI21X1_758/B vdd OAI21X1
XNOR2X1_273 INVX4_9/Y INVX1_140/A gnd NOR2X1_273/Y vdd NOR2X1
XNOR2X1_284 INVX1_57/A BUFX4_118/Y gnd NOR2X1_284/Y vdd NOR2X1
XOAI21X1_746 BUFX4_221/Y BUFX4_233/Y INVX2_128/A gnd OAI21X1_746/Y vdd OAI21X1
XOAI21X1_779 INVX2_132/Y BUFX4_85/Y OAI21X1_787/C gnd AOI21X1_266/B vdd OAI21X1
XOAI21X1_768 BUFX4_96/Y INVX8_18/Y AND2X2_31/A gnd NOR2X1_337/B vdd OAI21X1
XBUFX4_20 BUFX4_19/A gnd BUFX4_20/Y vdd BUFX4
XFILL_34_0_1 gnd vdd FILL
XBUFX4_86 wb_sel_i[0] gnd BUFX4_86/Y vdd BUFX4
XBUFX4_75 BUFX4_78/A gnd INVX8_1/A vdd BUFX4
XBUFX4_42 BUFX4_45/A gnd BUFX4_42/Y vdd BUFX4
XBUFX4_31 BUFX4_32/A gnd BUFX4_31/Y vdd BUFX4
XBUFX4_53 BUFX4_52/A gnd BUFX4_53/Y vdd BUFX4
XBUFX4_97 BUFX4_98/A gnd BUFX4_97/Y vdd BUFX4
XBUFX4_64 BUFX4_61/A gnd BUFX4_64/Y vdd BUFX4
XOR2X2_12 OR2X2_12/A OR2X2_12/B gnd OR2X2_12/Y vdd OR2X2
XOR2X2_5 OR2X2_5/A OR2X2_5/B gnd OR2X2_5/Y vdd OR2X2
XXNOR2X1_7 OR2X2_8/A BUFX4_112/Y gnd OR2X2_10/A vdd XNOR2X1
XFILL_25_0_1 gnd vdd FILL
XINVX8_12 BUFX4_35/Y gnd INVX8_12/Y vdd INVX8
XFILL_0_0_1 gnd vdd FILL
XINVX8_23 INVX8_23/A gnd OR2X2_18/B vdd INVX8
XOAI21X1_587 INVX2_54/Y BUFX4_161/Y OAI21X1_587/C gnd OAI21X1_588/B vdd OAI21X1
XOAI21X1_598 NOR2X1_280/Y INVX2_78/Y BUFX4_122/Y gnd AOI21X1_210/C vdd OAI21X1
XOAI21X1_554 AND2X2_27/Y INVX2_106/Y BUFX4_171/Y gnd OAI21X1_554/Y vdd OAI21X1
XOAI21X1_543 BUFX4_211/Y BUFX4_28/Y INVX2_73/A gnd OAI21X1_543/Y vdd OAI21X1
XOAI21X1_532 OAI21X1_532/A OAI21X1_532/B OAI21X1_528/Y gnd DFFSR_185/D vdd OAI21X1
XOAI21X1_576 NOR2X1_272/Y MUX2X1_1/B BUFX4_123/Y gnd AOI21X1_198/C vdd OAI21X1
XOAI21X1_565 INVX2_82/Y MUX2X1_6/S OAI21X1_333/C gnd AOI21X1_194/B vdd OAI21X1
XINVX1_7 INVX1_7/A gnd INVX1_7/Y vdd INVX1
XOAI21X1_510 BUFX4_57/Y NAND2X1_256/Y OAI21X1_510/C gnd AOI21X1_179/B vdd OAI21X1
XOAI21X1_521 BUFX4_167/Y OAI21X1_521/B BUFX4_38/Y gnd OAI21X1_522/B vdd OAI21X1
XFILL_8_1_1 gnd vdd FILL
XFILL_16_0_1 gnd vdd FILL
XOAI21X1_373 BUFX4_52/Y OAI21X1_373/B BUFX4_244/Y gnd OAI21X1_373/Y vdd OAI21X1
XOAI21X1_362 NOR2X1_212/Y INVX2_162/Y BUFX4_51/Y gnd OAI21X1_362/Y vdd OAI21X1
XAND2X2_7 AND2X2_7/A AND2X2_7/B gnd AND2X2_7/Y vdd AND2X2
XOAI21X1_340 AOI21X1_107/Y OAI21X1_339/Y OAI21X1_336/Y gnd DFFSR_239/D vdd OAI21X1
XOAI21X1_351 BUFX4_223/Y BUFX4_234/Y INVX2_165/A gnd OAI21X1_355/C vdd OAI21X1
XOAI21X1_384 BUFX4_222/Y BUFX4_233/Y INVX1_59/A gnd OAI21X1_384/Y vdd OAI21X1
XOAI21X1_395 INVX2_111/Y BUFX4_10/Y OAI21X1_621/C gnd OAI21X1_395/Y vdd OAI21X1
XAOI22X1_2 BUFX4_26/Y INVX1_9/A AOI22X1_2/C INVX8_6/Y gnd AOI22X1_2/Y vdd AOI22X1
XOAI21X1_192 INVX2_43/A INVX4_2/Y INVX1_85/A gnd AND2X2_10/A vdd OAI21X1
XOAI21X1_181 INVX4_11/A DFFSR_43/Q NAND2X1_103/Y gnd NOR2X1_51/A vdd OAI21X1
XOAI21X1_170 AND2X2_7/Y BUFX4_4/Y NAND2X1_95/Y gnd DFFSR_106/D vdd OAI21X1
XNAND2X1_12 BUFX4_165/Y wb_dat_i[19] gnd NAND2X1_12/Y vdd NAND2X1
XNAND2X1_67 DFFSR_139/Q AOI21X1_2/B gnd NAND2X1_67/Y vdd NAND2X1
XNAND2X1_45 AOI21X1_7/Y NOR2X1_10/Y gnd DFFSR_71/D vdd NAND2X1
XNAND2X1_34 wb_adr_i[4] wb_adr_i[3] gnd NAND2X1_34/Y vdd NAND2X1
XNAND2X1_56 NAND2X1_56/A NOR2X1_16/Y gnd DFFSR_77/D vdd NAND2X1
XNAND2X1_78 AND2X2_8/B NOR2X1_24/Y gnd OR2X2_4/A vdd NAND2X1
XNAND2X1_89 INVX1_70/Y AND2X2_5/B gnd AND2X2_6/A vdd NAND2X1
XNAND2X1_23 BUFX4_9/Y wb_dat_i[14] gnd OAI21X1_45/C vdd NAND2X1
XFILL_33_6_0 gnd vdd FILL
XAOI21X1_205 BUFX4_31/Y AOI21X1_205/B BUFX4_203/Y gnd AOI21X1_206/A vdd AOI21X1
XAOI21X1_216 INVX2_154/Y AOI21X1_216/B BUFX4_34/Y gnd OAI21X1_614/C vdd AOI21X1
XAOI22X1_10 BUFX4_25/Y INVX1_13/A INVX2_89/A INVX8_6/Y gnd NAND3X1_90/C vdd AOI22X1
XAOI21X1_238 BUFX4_32/Y AOI21X1_238/B BUFX4_206/Y gnd AOI21X1_239/A vdd AOI21X1
XAOI22X1_43 AOI22X1_43/A AOI21X1_61/Y AOI22X1_43/C AOI22X1_43/D gnd AOI22X1_43/Y vdd
+ AOI22X1
XAOI22X1_54 NOR2X1_190/Y AOI22X1_54/B AOI22X1_54/C NOR2X1_191/Y gnd AOI21X1_85/B vdd
+ AOI22X1
XAOI22X1_32 BUFX4_21/Y INVX1_8/A DFFSR_243/Q INVX8_6/Y gnd AOI22X1_32/Y vdd AOI22X1
XAOI22X1_21 BUFX4_21/Y INVX1_3/A INVX2_69/A INVX8_5/Y gnd NAND3X1_96/C vdd AOI22X1
XAOI21X1_249 NOR2X1_325/Y BUFX4_57/Y AOI21X1_249/C gnd OAI21X1_740/A vdd AOI21X1
XAOI22X1_76 INVX2_67/A INVX8_14/A INVX8_23/A INVX1_94/A gnd AOI22X1_76/Y vdd AOI22X1
XAOI22X1_65 INVX1_54/A INVX8_17/A INVX8_23/A INVX1_97/A gnd AOI22X1_65/Y vdd AOI22X1
XAOI21X1_227 INVX2_97/Y OAI21X1_628/B BUFX4_34/Y gnd AOI21X1_227/Y vdd AOI21X1
XFILL_24_6_0 gnd vdd FILL
XNAND3X1_209 OAI21X1_314/Y OAI21X1_315/Y AOI22X1_68/Y gnd AOI22X1_77/C vdd NAND3X1
XOAI22X1_5 BUFX4_78/Y INVX2_11/Y INVX1_30/Y OAI22X1_1/D gnd NOR2X1_6/A vdd OAI22X1
XFILL_15_6_0 gnd vdd FILL
XDFFSR_229 AOI22X1_4/C CLKBUF1_6/Y BUFX4_130/Y vdd DFFSR_229/D gnd vdd DFFSR
XDFFSR_218 INVX1_43/A DFFSR_8/CLK DFFSR_151/R vdd DFFSR_218/D gnd vdd DFFSR
XDFFSR_207 INVX2_110/A CLKBUF1_26/Y DFFSR_194/R vdd DFFSR_207/D gnd vdd DFFSR
XINVX2_14 DFFSR_6/Q gnd INVX2_14/Y vdd INVX2
XINVX2_36 INVX2_36/A gnd INVX2_36/Y vdd INVX2
XINVX2_58 INVX1_41/A gnd INVX2_58/Y vdd INVX2
XINVX2_47 INVX2_47/A gnd INVX2_47/Y vdd INVX2
XINVX2_69 INVX2_69/A gnd INVX2_69/Y vdd INVX2
XINVX2_25 DFFSR_57/Q gnd INVX2_25/Y vdd INVX2
XFILL_30_4_0 gnd vdd FILL
XNAND2X1_219 BUFX4_165/Y wb_dat_i[20] gnd NAND2X1_219/Y vdd NAND2X1
XNAND2X1_208 BUFX4_73/Y wb_dat_i[26] gnd OAI21X1_572/C vdd NAND2X1
XBUFX4_181 AND2X2_1/Y gnd BUFX4_181/Y vdd BUFX4
XNOR2X1_263 INVX4_8/Y INVX1_136/Y gnd NOR2X1_263/Y vdd NOR2X1
XNOR2X1_252 INVX4_7/Y INVX1_137/Y gnd NOR2X1_252/Y vdd NOR2X1
XNOR2X1_274 INVX4_9/Y OR2X2_17/A gnd NOR2X1_274/Y vdd NOR2X1
XNOR2X1_230 INVX1_28/A BUFX4_241/Y gnd NOR2X1_230/Y vdd NOR2X1
XBUFX4_170 INVX8_19/Y gnd BUFX4_170/Y vdd BUFX4
XNOR2X1_285 INVX1_52/A BUFX4_118/Y gnd NOR2X1_285/Y vdd NOR2X1
XNOR2X1_241 BUFX4_148/Y NOR2X1_224/A gnd INVX1_134/A vdd NOR2X1
XBUFX4_192 BUFX4_193/A gnd BUFX4_192/Y vdd BUFX4
XOAI21X1_714 OAI21X1_714/A BUFX4_208/Y OAI21X1_714/C gnd DFFSR_122/D vdd OAI21X1
XFILL_21_4_0 gnd vdd FILL
XOAI21X1_725 NOR2X1_321/Y OAI21X1_725/B OAI21X1_725/C gnd DFFSR_119/D vdd OAI21X1
XOAI21X1_747 NOR2X1_327/Y INVX2_128/Y BUFX4_51/Y gnd AOI21X1_251/C vdd OAI21X1
XNOR2X1_296 INVX8_22/Y NOR2X1_296/B gnd INVX1_141/A vdd NOR2X1
XOAI21X1_758 BUFX4_167/Y OAI21X1_758/B BUFX4_38/Y gnd OAI21X1_759/B vdd OAI21X1
XOAI21X1_736 BUFX4_99/Y INVX4_6/Y INVX1_112/A gnd NOR2X1_329/B vdd OAI21X1
XOAI21X1_769 BUFX4_62/Y AOI21X1_258/B OAI21X1_769/C gnd AOI21X1_260/B vdd OAI21X1
XOAI21X1_703 INVX1_146/Y OR2X2_18/B MUX2X1_2/A gnd OAI21X1_704/C vdd OAI21X1
XFILL_29_5_0 gnd vdd FILL
XFILL_4_5_0 gnd vdd FILL
XINVX8_1 INVX8_1/A gnd INVX8_1/Y vdd INVX8
XFILL_12_4_0 gnd vdd FILL
XBUFX4_32 BUFX4_32/A gnd BUFX4_32/Y vdd BUFX4
XBUFX4_10 wb_sel_i[1] gnd BUFX4_10/Y vdd BUFX4
XBUFX4_21 INVX8_1/Y gnd BUFX4_21/Y vdd BUFX4
XBUFX4_43 BUFX4_45/A gnd BUFX4_43/Y vdd BUFX4
XBUFX4_98 BUFX4_98/A gnd BUFX4_98/Y vdd BUFX4
XBUFX4_76 BUFX4_78/A gnd BUFX4_76/Y vdd BUFX4
XBUFX4_65 BUFX4_61/A gnd BUFX4_65/Y vdd BUFX4
XBUFX4_87 INVX8_8/Y gnd BUFX4_87/Y vdd BUFX4
XBUFX4_54 BUFX4_52/A gnd BUFX4_54/Y vdd BUFX4
XXNOR2X1_8 XNOR2X1_8/A INVX2_43/Y gnd XNOR2X1_8/Y vdd XNOR2X1
XOR2X2_13 OR2X2_12/A OR2X2_13/B gnd OR2X2_13/Y vdd OR2X2
XOR2X2_6 OR2X2_6/A OR2X2_6/B gnd OR2X2_6/Y vdd OR2X2
XINVX8_13 INVX8_13/A gnd INVX8_13/Y vdd INVX8
XINVX8_24 wb_rst_i gnd INVX8_24/Y vdd INVX8
XOAI21X1_588 BUFX4_121/Y OAI21X1_588/B BUFX4_114/Y gnd OAI21X1_589/B vdd OAI21X1
XOAI21X1_599 INVX2_78/Y BUFX4_165/Y NAND2X1_224/Y gnd OAI21X1_599/Y vdd OAI21X1
XOAI21X1_555 INVX2_106/Y BUFX4_83/Y OAI21X1_732/C gnd OAI21X1_556/B vdd OAI21X1
XOAI21X1_544 NOR2X1_263/Y INVX2_73/Y BUFX4_170/Y gnd AOI21X1_186/C vdd OAI21X1
XOAI21X1_533 INVX8_21/A BUFX4_33/Y INVX1_36/A gnd OAI21X1_533/Y vdd OAI21X1
XOAI21X1_577 MUX2X1_1/B BUFX4_70/Y OAI21X1_458/C gnd OAI21X1_577/Y vdd OAI21X1
XOAI21X1_566 AND2X2_29/Y INVX2_109/Y BUFX4_119/Y gnd AOI21X1_196/C vdd OAI21X1
XINVX1_8 INVX1_8/A gnd INVX1_8/Y vdd INVX1
XOAI21X1_511 INVX2_72/Y BUFX4_5/Y NAND2X1_236/Y gnd OAI21X1_512/B vdd OAI21X1
XOAI21X1_522 OAI21X1_522/A OAI21X1_522/B OAI21X1_522/C gnd DFFSR_188/D vdd OAI21X1
XOAI21X1_500 BUFX4_166/Y OAI21X1_500/B BUFX4_39/Y gnd OAI21X1_501/B vdd OAI21X1
XFILL_9_1 gnd vdd FILL
XFILL_35_3_0 gnd vdd FILL
XFILL_26_3_0 gnd vdd FILL
XFILL_1_3_0 gnd vdd FILL
XOAI21X1_330 OAI21X1_330/A OAI21X1_329/Y OAI21X1_330/C gnd DFFSR_241/D vdd OAI21X1
XOAI21X1_341 BUFX4_224/Y BUFX4_231/Y INVX2_67/A gnd OAI21X1_341/Y vdd OAI21X1
XOAI21X1_374 OAI21X1_374/A OAI21X1_373/Y OAI21X1_374/C gnd DFFSR_230/D vdd OAI21X1
XOAI21X1_363 INVX2_162/Y BUFX4_164/Y NAND2X1_216/Y gnd OAI21X1_364/B vdd OAI21X1
XOAI21X1_396 BUFX4_223/Y BUFX4_234/Y INVX1_50/A gnd OAI21X1_400/C vdd OAI21X1
XOAI21X1_352 NOR2X1_210/Y INVX2_165/Y BUFX4_56/Y gnd OAI21X1_352/Y vdd OAI21X1
XAND2X2_8 AND2X2_8/A AND2X2_8/B gnd AND2X2_8/Y vdd AND2X2
XOAI21X1_385 NOR2X1_219/Y INVX2_153/Y BUFX4_56/Y gnd AOI21X1_127/C vdd OAI21X1
XFILL_9_4_0 gnd vdd FILL
XFILL_17_3_0 gnd vdd FILL
XAOI22X1_3 DFFSR_165/Q AOI22X1_1/B INVX8_5/Y AOI22X1_3/D gnd AOI22X1_3/Y vdd AOI22X1
XOAI21X1_182 INVX8_9/Y DFFSR_33/Q INVX2_44/Y gnd OAI21X1_183/C vdd OAI21X1
XOAI21X1_160 OR2X2_4/Y NAND2X1_86/Y BUFX4_97/Y gnd BUFX4_1/A vdd OAI21X1
XOAI21X1_171 AOI21X1_22/Y BUFX4_4/Y NAND2X1_96/Y gnd DFFSR_107/D vdd OAI21X1
XOAI21X1_193 AND2X2_10/Y NOR2X1_59/Y BUFX4_248/Y gnd OAI21X1_194/C vdd OAI21X1
XNAND2X1_13 BUFX4_160/Y wb_dat_i[20] gnd NAND2X1_13/Y vdd NAND2X1
XNAND2X1_46 NAND2X1_46/A NAND2X1_46/B gnd AOI21X1_8/C vdd NAND2X1
XNAND2X1_35 INVX2_39/Y NOR2X1_3/Y gnd NOR2X1_19/B vdd NAND2X1
XNAND2X1_57 NAND2X1_57/A NOR2X1_17/Y gnd DFFSR_78/D vdd NAND2X1
XNAND2X1_68 INVX1_120/A BUFX4_190/Y gnd NAND3X1_94/B vdd NAND2X1
XNAND2X1_79 INVX1_78/A NOR2X1_26/Y gnd OR2X2_4/B vdd NAND2X1
XNAND2X1_24 BUFX4_11/Y wb_dat_i[15] gnd OAI21X1_47/C vdd NAND2X1
XFILL_33_6_1 gnd vdd FILL
XFILL_32_1_0 gnd vdd FILL
XAOI21X1_239 AOI21X1_239/A OAI21X1_638/Y NOR2X1_292/Y gnd DFFSR_151/D vdd AOI21X1
XAOI21X1_228 BUFX4_31/Y AOI21X1_228/B BUFX4_203/Y gnd AOI21X1_229/A vdd AOI21X1
XAOI21X1_206 AOI21X1_206/A AOI21X1_206/B NOR2X1_277/Y gnd DFFSR_168/D vdd AOI21X1
XAOI21X1_217 BUFX4_34/Y AOI21X1_217/B BUFX4_210/Y gnd AOI21X1_218/A vdd AOI21X1
XAOI22X1_66 AOI21X1_94/Y AOI22X1_66/B AOI22X1_66/C AOI22X1_66/D gnd AOI22X1_66/Y vdd
+ AOI22X1
XAOI22X1_11 INVX8_6/Y DFFSR_233/Q INVX2_160/A INVX8_5/Y gnd AOI22X1_11/Y vdd AOI22X1
XNOR3X1_1 wb_adr_i[4] wb_adr_i[3] INVX4_1/Y gnd NOR3X1_1/Y vdd NOR3X1
XAOI22X1_55 AOI21X1_86/Y AOI22X1_55/B AOI22X1_55/C AOI22X1_55/D gnd AOI22X1_55/Y vdd
+ AOI22X1
XAOI22X1_22 INVX2_68/A BUFX4_124/Y INVX8_6/Y INVX2_67/A gnd NAND3X1_96/A vdd AOI22X1
XAOI22X1_33 INVX1_69/Y BUFX4_2/Y OR2X2_5/Y AOI21X1_24/Y gnd DFFSR_111/D vdd AOI22X1
XAOI22X1_77 AOI22X1_77/A INVX1_111/A AOI22X1_77/C INVX1_122/A gnd AOI22X1_77/Y vdd
+ AOI22X1
XAOI22X1_44 AOI22X1_44/A AOI21X1_63/Y AOI21X1_64/Y AOI22X1_44/D gnd AOI22X1_44/Y vdd
+ AOI22X1
XFILL_24_6_1 gnd vdd FILL
XFILL_23_1_0 gnd vdd FILL
XOAI22X1_6 OAI22X1_4/A INVX2_33/Y OAI22X1_4/C INVX1_31/Y gnd NOR2X1_6/B vdd OAI22X1
XFILL_6_2_0 gnd vdd FILL
XFILL_15_6_1 gnd vdd FILL
XFILL_14_1_0 gnd vdd FILL
XDFFSR_219 INVX1_44/A CLKBUF1_37/Y DFFSR_198/R vdd DFFSR_219/D gnd vdd DFFSR
XDFFSR_208 INVX2_83/A CLKBUF1_24/Y DFFSR_194/R vdd DFFSR_208/D gnd vdd DFFSR
XINVX2_15 DFFSR_7/Q gnd INVX2_15/Y vdd INVX2
XINVX2_26 INVX2_26/A gnd INVX2_26/Y vdd INVX2
XINVX2_48 INVX2_48/A gnd INVX2_48/Y vdd INVX2
XINVX2_37 INVX2_37/A gnd INVX2_37/Y vdd INVX2
XINVX2_59 INVX1_42/A gnd INVX2_59/Y vdd INVX2
XFILL_30_4_1 gnd vdd FILL
XNAND2X1_209 INVX1_125/Y NOR2X1_191/Y gnd NOR2X1_239/B vdd NAND2X1
XBUFX4_160 wb_sel_i[2] gnd BUFX4_160/Y vdd BUFX4
XBUFX4_193 BUFX4_193/A gnd AOI21X1_1/B vdd BUFX4
XNOR2X1_275 DFFSR_169/Q BUFX4_114/Y gnd NOR2X1_275/Y vdd NOR2X1
XNOR2X1_264 INVX4_8/Y INVX1_137/Y gnd NOR2X1_264/Y vdd NOR2X1
XNOR2X1_231 INVX1_26/A BUFX4_241/Y gnd NOR2X1_231/Y vdd NOR2X1
XBUFX4_171 INVX8_19/Y gnd BUFX4_171/Y vdd BUFX4
XNOR2X1_253 BUFX4_152/Y INVX1_129/A gnd AND2X2_27/A vdd NOR2X1
XBUFX4_182 AND2X2_1/Y gnd BUFX4_182/Y vdd BUFX4
XNOR2X1_297 INVX1_141/Y BUFX4_63/Y gnd NOR2X1_297/Y vdd NOR2X1
XNOR2X1_286 INVX1_51/A BUFX4_117/Y gnd NOR2X1_286/Y vdd NOR2X1
XNOR2X1_242 INVX4_7/Y INVX1_134/Y gnd NOR2X1_242/Y vdd NOR2X1
XNOR2X1_220 OR2X2_12/A INVX1_124/Y gnd NOR2X1_220/Y vdd NOR2X1
XOAI21X1_715 INVX1_102/Y BUFX4_84/Y NAND2X1_240/Y gnd OAI21X1_715/Y vdd OAI21X1
XOAI21X1_726 INVX2_74/Y BUFX4_79/Y NAND2X1_244/Y gnd NAND2X1_322/B vdd OAI21X1
XFILL_21_4_1 gnd vdd FILL
XOAI21X1_748 INVX2_128/Y BUFX4_162/Y NAND2X1_330/Y gnd OAI21X1_749/B vdd OAI21X1
XOAI21X1_737 NOR2X1_325/Y INVX2_127/Y BUFX4_168/Y gnd AOI21X1_249/C vdd OAI21X1
XOAI21X1_759 OAI21X1_759/A OAI21X1_759/B OAI21X1_755/Y gnd DFFSR_195/D vdd OAI21X1
XOAI21X1_704 BUFX4_64/Y OAI21X1_704/B OAI21X1_704/C gnd OAI21X1_706/A vdd OAI21X1
XFILL_29_5_1 gnd vdd FILL
XFILL_28_0_0 gnd vdd FILL
XFILL_3_0_0 gnd vdd FILL
XFILL_4_5_1 gnd vdd FILL
XINVX8_2 INVX8_2/A gnd INVX8_2/Y vdd INVX8
XFILL_12_4_1 gnd vdd FILL
XBUFX4_33 BUFX4_32/A gnd BUFX4_33/Y vdd BUFX4
XBUFX4_66 BUFX4_61/A gnd BUFX4_66/Y vdd BUFX4
XBUFX4_77 BUFX4_78/A gnd BUFX4_77/Y vdd BUFX4
XBUFX4_11 wb_sel_i[1] gnd BUFX4_11/Y vdd BUFX4
XBUFX4_22 INVX8_1/Y gnd BUFX4_22/Y vdd BUFX4
XBUFX4_44 BUFX4_45/A gnd BUFX4_44/Y vdd BUFX4
XBUFX4_55 BUFX4_52/A gnd BUFX4_55/Y vdd BUFX4
XFILL_19_0_0 gnd vdd FILL
XBUFX4_88 INVX8_8/Y gnd DFFSR_98/R vdd BUFX4
XBUFX4_99 BUFX4_98/A gnd BUFX4_99/Y vdd BUFX4
XOR2X2_14 OR2X2_14/A INVX4_7/Y gnd OR2X2_14/Y vdd OR2X2
XOR2X2_7 OR2X2_7/A OR2X2_7/B gnd OR2X2_7/Y vdd OR2X2
XINVX2_160 INVX2_160/A gnd INVX2_160/Y vdd INVX2
XXNOR2X1_9 XNOR2X1_9/A OR2X2_9/B gnd INVX1_105/A vdd XNOR2X1
XINVX1_9 INVX1_9/A gnd INVX1_9/Y vdd INVX1
XOAI21X1_523 BUFX4_206/Y BUFX4_32/Y INVX1_42/A gnd OAI21X1_523/Y vdd OAI21X1
XINVX8_14 INVX8_14/A gnd INVX8_14/Y vdd INVX8
XOAI21X1_512 BUFX4_222/Y OAI21X1_512/B BUFX4_49/Y gnd AOI21X1_179/A vdd OAI21X1
XOAI21X1_501 AOI21X1_174/Y OAI21X1_501/B OAI21X1_497/Y gnd DFFSR_193/D vdd OAI21X1
XOAI21X1_589 OAI21X1_589/A OAI21X1_589/B NAND2X1_264/Y gnd DFFSR_170/D vdd OAI21X1
XOAI21X1_556 BUFX4_171/Y OAI21X1_556/B BUFX4_36/Y gnd OAI21X1_557/B vdd OAI21X1
XOAI21X1_545 INVX2_73/Y BUFX4_81/Y NAND2X1_244/Y gnd OAI21X1_546/B vdd OAI21X1
XOAI21X1_534 NOR2X1_261/Y INVX2_95/Y BUFX4_166/Y gnd AOI21X1_184/C vdd OAI21X1
XOAI21X1_578 BUFX4_123/Y OAI21X1_577/Y BUFX4_116/Y gnd OAI21X1_578/Y vdd OAI21X1
XOAI21X1_567 INVX2_109/Y MUX2X1_7/S OAI21X1_567/C gnd OAI21X1_568/B vdd OAI21X1
XFILL_9_2 gnd vdd FILL
XFILL_35_3_1 gnd vdd FILL
XNAND3X1_190 OAI21X1_277/Y XNOR2X1_10/Y INVX1_108/A gnd AOI21X1_45/B vdd NAND3X1
XFILL_26_3_1 gnd vdd FILL
XFILL_1_3_1 gnd vdd FILL
XOAI21X1_364 BUFX4_51/Y OAI21X1_364/B BUFX4_243/Y gnd OAI21X1_365/B vdd OAI21X1
XOAI21X1_331 BUFX4_224/Y BUFX4_231/Y INVX2_81/A gnd OAI21X1_331/Y vdd OAI21X1
XOAI21X1_320 OAI21X1_320/A OAI21X1_319/Y OAI21X1_267/Y gnd DFFSR_243/D vdd OAI21X1
XOAI21X1_342 NOR2X1_208/Y INVX2_67/Y BUFX4_55/Y gnd AOI21X1_108/C vdd OAI21X1
XOAI21X1_353 INVX2_165/Y BUFX4_71/Y OAI21X1_353/C gnd OAI21X1_354/B vdd OAI21X1
XAND2X2_9 OR2X2_8/A OR2X2_8/B gnd AND2X2_9/Y vdd AND2X2
XOAI21X1_375 BUFX4_220/Y BUFX4_230/Y AOI22X1_4/C gnd OAI21X1_379/C vdd OAI21X1
XOAI21X1_397 NOR2X1_222/Y INVX2_70/Y BUFX4_56/Y gnd AOI21X1_132/C vdd OAI21X1
XFILL_9_4_1 gnd vdd FILL
XOAI21X1_386 INVX2_153/Y BUFX4_6/Y NAND2X1_232/Y gnd OAI21X1_387/B vdd OAI21X1
XFILL_17_3_1 gnd vdd FILL
XOAI21X1_150 BUFX4_93/Y BUFX4_103/Y INVX1_16/A gnd BUFX2_26/A vdd OAI21X1
XOAI21X1_194 INVX2_18/A INVX1_107/A OAI21X1_194/C gnd INVX4_4/A vdd OAI21X1
XAOI22X1_4 BUFX4_25/Y INVX1_10/A AOI22X1_4/C INVX8_6/Y gnd AOI22X1_4/Y vdd AOI22X1
XOAI21X1_183 INVX1_81/Y INVX8_9/Y OAI21X1_183/C gnd INVX1_82/A vdd OAI21X1
XOAI21X1_172 NOR2X1_43/Y AND2X2_8/A NOR2X1_46/B gnd OAI21X1_173/C vdd OAI21X1
XOAI21X1_161 XOR2X1_1/A BUFX4_3/Y NAND2X1_87/Y gnd DFFSR_100/D vdd OAI21X1
XNAND2X1_14 BUFX4_162/Y wb_dat_i[21] gnd OAI21X1_27/C vdd NAND2X1
XNAND2X1_25 wb_dat_i[0] BUFX4_79/Y gnd NAND2X1_25/Y vdd NAND2X1
XNAND2X1_36 NAND3X1_69/Y NAND3X1_70/Y gnd AOI21X1_1/C vdd NAND2X1
XNAND2X1_47 AOI21X1_8/Y NOR2X1_11/Y gnd DFFSR_72/D vdd NAND2X1
XNAND2X1_69 DFFSR_141/Q BUFX4_192/Y gnd NAND3X1_95/A vdd NAND2X1
XNAND2X1_58 AOI21X1_16/Y NAND2X1_58/B gnd DFFSR_79/D vdd NAND2X1
XFILL_32_1_1 gnd vdd FILL
XAOI22X1_12 DFFSR_169/Q AOI22X1_1/B BUFX4_25/Y DFFSR_22/Q gnd AOI22X1_12/Y vdd AOI22X1
XAOI21X1_207 INVX2_121/Y NAND2X1_266/Y BUFX4_31/Y gnd OAI21X1_595/C vdd AOI21X1
XAOI21X1_229 AOI21X1_229/A OAI21X1_628/Y NOR2X1_288/Y gnd DFFSR_156/D vdd AOI21X1
XAOI22X1_23 INVX2_109/A BUFX4_124/Y INVX8_5/Y INVX2_110/A gnd NAND3X1_97/B vdd AOI22X1
XAOI21X1_218 AOI21X1_218/A AOI21X1_218/B NOR2X1_284/Y gnd DFFSR_161/D vdd AOI21X1
XAOI22X1_67 AOI21X1_98/Y AOI22X1_67/B AOI22X1_67/C AOI21X1_99/Y gnd AOI22X1_67/Y vdd
+ AOI22X1
XAOI22X1_56 AOI22X1_56/A AOI22X1_56/B AOI22X1_56/C AOI22X1_56/D gnd AOI22X1_56/Y vdd
+ AOI22X1
XAOI22X1_78 BUFX4_207/Y MUX2X1_5/Y AOI22X1_78/C AOI22X1_78/D gnd DFFSR_145/D vdd AOI22X1
XNOR3X1_2 NOR3X1_2/A NOR3X1_2/B NOR3X1_2/C gnd AND2X2_8/A vdd NOR3X1
XAOI22X1_34 INVX1_66/Y BUFX4_2/Y NOR2X1_45/Y AOI22X1_34/D gnd DFFSR_112/D vdd AOI22X1
XAOI22X1_45 AOI22X1_45/A AOI21X1_65/Y AOI21X1_66/Y AOI22X1_45/D gnd AOI22X1_45/Y vdd
+ AOI22X1
XFILL_23_1_1 gnd vdd FILL
XOAI22X1_7 INVX8_1/A INVX2_12/Y INVX2_34/Y OAI22X1_7/D gnd NOR2X1_7/A vdd OAI22X1
XFILL_6_2_1 gnd vdd FILL
XFILL_14_1_1 gnd vdd FILL
XDFFSR_209 DFFSR_209/Q CLKBUF1_32/A DFFSR_236/R vdd DFFSR_209/D gnd vdd DFFSR
XINVX2_49 INVX2_49/A gnd INVX2_49/Y vdd INVX2
XINVX2_16 DFFSR_8/Q gnd INVX2_16/Y vdd INVX2
XINVX2_38 DFFSR_54/Q gnd INVX2_38/Y vdd INVX2
XINVX2_27 INVX2_27/A gnd INVX2_27/Y vdd INVX2
XCLKBUF1_1 CLKBUF1_5/A gnd CLKBUF1_1/Y vdd CLKBUF1
XBUFX4_161 wb_sel_i[2] gnd BUFX4_161/Y vdd BUFX4
XBUFX4_172 BUFX4_172/A gnd BUFX4_172/Y vdd BUFX4
XBUFX4_150 BUFX4_152/A gnd BUFX4_150/Y vdd BUFX4
XBUFX4_194 BUFX4_194/A gnd BUFX4_194/Y vdd BUFX4
XNOR2X1_254 DFFSR_196/Q BUFX4_36/Y gnd NOR2X1_254/Y vdd NOR2X1
XNOR2X1_243 BUFX4_152/Y NOR2X1_243/B gnd AND2X2_25/A vdd NOR2X1
XBUFX4_183 AND2X2_1/Y gnd BUFX4_183/Y vdd BUFX4
XNOR2X1_276 INVX8_19/A OR2X2_15/A gnd NOR2X1_276/Y vdd NOR2X1
XNOR2X1_232 INVX2_66/A BUFX4_35/Y gnd NOR2X1_232/Y vdd NOR2X1
XNOR2X1_298 INVX8_22/Y NOR2X1_316/B gnd INVX1_142/A vdd NOR2X1
XNOR2X1_265 BUFX4_231/Y INVX1_131/A gnd AND2X2_28/A vdd NOR2X1
XNOR2X1_221 INVX1_54/A BUFX4_240/Y gnd NOR2X1_221/Y vdd NOR2X1
XNOR2X1_210 NOR2X1_224/A INVX8_14/Y gnd NOR2X1_210/Y vdd NOR2X1
XOAI21X1_705 MUX2X1_2/A BUFX4_12/Y OAI21X1_515/C gnd NAND2X1_312/B vdd OAI21X1
XNOR2X1_287 OR2X2_17/B NOR2X1_287/B gnd NOR2X1_287/Y vdd NOR2X1
XOAI21X1_716 INVX1_158/Y DFFSR_121/Q BUFX4_113/Y gnd OAI21X1_716/Y vdd OAI21X1
XOAI21X1_727 INVX1_159/Y INVX2_74/A BUFX4_114/Y gnd OAI21X1_728/B vdd OAI21X1
XOAI21X1_738 INVX2_127/Y BUFX4_72/Y OAI21X1_738/C gnd OAI21X1_738/Y vdd OAI21X1
XOAI21X1_749 BUFX4_51/Y OAI21X1_749/B BUFX4_243/Y gnd OAI21X1_750/B vdd OAI21X1
XFILL_28_0_1 gnd vdd FILL
XFILL_3_0_1 gnd vdd FILL
XINVX8_3 INVX8_3/A gnd INVX8_3/Y vdd INVX8
XBUFX4_45 BUFX4_45/A gnd BUFX4_45/Y vdd BUFX4
XBUFX4_78 BUFX4_78/A gnd BUFX4_78/Y vdd BUFX4
XFILL_19_0_1 gnd vdd FILL
XBUFX4_23 INVX8_1/Y gnd BUFX4_23/Y vdd BUFX4
XBUFX4_56 BUFX4_52/A gnd BUFX4_56/Y vdd BUFX4
XBUFX4_89 INVX8_8/Y gnd BUFX4_89/Y vdd BUFX4
XBUFX4_34 BUFX4_32/A gnd BUFX4_34/Y vdd BUFX4
XBUFX4_67 BUFX4_61/A gnd BUFX4_67/Y vdd BUFX4
XBUFX4_12 wb_sel_i[1] gnd BUFX4_12/Y vdd BUFX4
XOR2X2_15 OR2X2_15/A INVX4_7/Y gnd OR2X2_15/Y vdd OR2X2
XINVX2_150 INVX2_150/A gnd INVX2_150/Y vdd INVX2
XOR2X2_8 OR2X2_8/A OR2X2_8/B gnd OR2X2_8/Y vdd OR2X2
XINVX2_161 DFFSR_137/Q gnd INVX2_161/Y vdd INVX2
XOAI21X1_557 AOI21X1_188/Y OAI21X1_557/B OAI21X1_553/Y gnd DFFSR_180/D vdd OAI21X1
XOAI21X1_546 BUFX4_171/Y OAI21X1_546/B BUFX4_36/Y gnd OAI21X1_547/B vdd OAI21X1
XOAI21X1_524 AND2X2_25/Y INVX2_59/Y BUFX4_169/Y gnd AOI21X1_182/C vdd OAI21X1
XOAI21X1_535 INVX2_95/Y BUFX4_79/Y NAND2X1_242/Y gnd OAI21X1_535/Y vdd OAI21X1
XINVX8_15 INVX8_15/A gnd BUFX4_52/A vdd INVX8
XOAI21X1_502 BUFX4_203/Y BUFX4_30/Y INVX2_86/A gnd OAI21X1_502/Y vdd OAI21X1
XOAI21X1_513 BUFX4_203/Y BUFX4_30/Y DFFSR_189/Q gnd OAI21X1_513/Y vdd OAI21X1
XOAI21X1_579 AOI21X1_198/Y OAI21X1_578/Y NAND2X1_262/Y gnd DFFSR_173/D vdd OAI21X1
XOAI21X1_568 BUFX4_119/Y OAI21X1_568/B BUFX4_116/Y gnd OAI21X1_569/B vdd OAI21X1
XFILL_9_3 gnd vdd FILL
XNAND3X1_180 INVX2_42/Y INVX8_13/A AOI21X1_36/B gnd NAND3X1_180/Y vdd NAND3X1
XNAND3X1_191 BUFX4_248/Y NAND3X1_191/B NAND3X1_191/C gnd NAND3X1_191/Y vdd NAND3X1
XOAI21X1_310 INVX2_79/A BUFX4_176/Y AOI21X1_96/Y gnd OAI21X1_310/Y vdd OAI21X1
XOAI21X1_376 NOR2X1_216/Y INVX2_148/Y BUFX4_52/Y gnd OAI21X1_376/Y vdd OAI21X1
XOAI21X1_365 OAI21X1_365/A OAI21X1_365/B OAI21X1_365/C gnd DFFSR_233/D vdd OAI21X1
XOAI21X1_321 BUFX4_223/Y BUFX4_234/Y INVX2_65/A gnd OAI21X1_325/C vdd OAI21X1
XOAI21X1_343 INVX2_67/Y MUX2X1_6/S OAI21X1_572/C gnd OAI21X1_343/Y vdd OAI21X1
XOAI21X1_354 BUFX4_53/Y OAI21X1_354/B BUFX4_242/Y gnd OAI21X1_354/Y vdd OAI21X1
XOAI21X1_398 INVX2_70/Y BUFX4_12/Y NAND2X1_236/Y gnd OAI21X1_399/B vdd OAI21X1
XOAI21X1_332 NOR2X1_206/Y INVX2_81/Y BUFX4_56/Y gnd AOI21X1_106/C vdd OAI21X1
XOAI21X1_387 BUFX4_54/Y OAI21X1_387/B BUFX4_242/Y gnd OAI21X1_388/B vdd OAI21X1
XFILL_27_6_0 gnd vdd FILL
XFILL_2_6_0 gnd vdd FILL
XOAI21X1_195 NOR2X1_48/B INVX2_48/A INVX2_42/A gnd AOI21X1_46/A vdd OAI21X1
XAOI22X1_5 BUFX4_25/Y INVX1_11/A INVX2_79/A INVX8_5/Y gnd AOI22X1_5/Y vdd AOI22X1
XOAI21X1_184 INVX2_44/Y DFFSR_33/Q XNOR2X1_3/Y gnd INVX1_83/A vdd OAI21X1
XOAI21X1_140 BUFX4_95/Y BUFX4_102/Y INVX2_6/A gnd BUFX2_16/A vdd OAI21X1
XOAI21X1_151 BUFX4_94/Y BUFX4_97/Y INVX1_1/A gnd BUFX2_27/A vdd OAI21X1
XOAI21X1_173 INVX1_73/Y NOR2X1_46/B OAI21X1_173/C gnd DFFSR_108/D vdd OAI21X1
XFILL_10_5_0 gnd vdd FILL
XOAI21X1_162 BUFX4_3/Y XOR2X1_1/Y NAND2X1_88/Y gnd DFFSR_101/D vdd OAI21X1
XNAND2X1_15 BUFX4_164/Y wb_dat_i[22] gnd OAI21X1_29/C vdd NAND2X1
XNAND2X1_37 AOI21X1_1/Y NOR2X1_2/Y gnd DFFSR_65/D vdd NAND2X1
XNAND2X1_26 BUFX4_81/Y wb_dat_i[1] gnd NAND2X1_26/Y vdd NAND2X1
XNAND2X1_48 NAND3X1_78/Y NAND2X1_48/B gnd AOI21X1_9/C vdd NAND2X1
XNAND2X1_59 NAND2X1_59/A NAND2X1_59/B gnd DFFSR_80/D vdd NAND2X1
XFILL_18_6_0 gnd vdd FILL
XNAND2X1_190 AOI22X1_60/Y AOI22X1_61/Y gnd NAND2X1_190/Y vdd NAND2X1
XAOI22X1_13 INVX2_54/A AOI22X1_7/B INVX8_5/Y INVX2_55/A gnd NAND3X1_92/B vdd AOI22X1
XAOI22X1_57 AOI22X1_57/A NOR2X1_189/Y NOR2X1_190/Y AOI22X1_57/D gnd AOI22X1_57/Y vdd
+ AOI22X1
XAOI21X1_208 BUFX4_31/Y OAI21X1_596/Y BUFX4_203/Y gnd AOI21X1_209/A vdd AOI21X1
XAOI22X1_46 AOI22X1_46/A NOR2X1_190/Y NOR2X1_191/Y AOI22X1_46/D gnd AOI22X1_46/Y vdd
+ AOI22X1
XAOI22X1_24 BUFX4_21/Y INVX1_4/A DFFSR_239/Q INVX8_6/Y gnd NAND3X1_97/C vdd AOI22X1
XAOI22X1_35 INVX1_67/Y BUFX4_4/Y OR2X2_6/Y AOI22X1_35/D gnd DFFSR_113/D vdd AOI22X1
XAOI21X1_219 AND2X2_30/Y BUFX4_57/Y AOI21X1_219/C gnd OAI21X1_619/A vdd AOI21X1
XAOI22X1_68 AOI22X1_68/A NOR2X1_189/Y NOR2X1_190/Y AOI22X1_68/D gnd AOI22X1_68/Y vdd
+ AOI22X1
XAOI22X1_79 BUFX4_212/Y MUX2X1_6/Y AOI22X1_79/C AOI22X1_79/D gnd DFFSR_144/D vdd AOI22X1
XNOR3X1_3 NOR3X1_3/A NOR3X1_3/B NOR3X1_3/C gnd NOR3X1_3/Y vdd NOR3X1
XOAI22X1_8 OAI22X1_4/C INVX1_32/Y INVX1_33/Y INVX8_5/A gnd NOR2X1_7/B vdd OAI22X1
XAOI21X1_90 INVX2_128/Y BUFX4_156/Y AOI21X1_71/C gnd AOI22X1_56/A vdd AOI21X1
XFILL_33_4_0 gnd vdd FILL
XFILL_19_1 gnd vdd FILL
XINVX2_17 wb_adr_i[3] gnd INVX2_17/Y vdd INVX2
XINVX2_39 wb_adr_i[4] gnd INVX2_39/Y vdd INVX2
XINVX2_28 INVX2_28/A gnd INVX2_28/Y vdd INVX2
XFILL_24_4_0 gnd vdd FILL
XFILL_7_5_0 gnd vdd FILL
XFILL_15_4_0 gnd vdd FILL
XMUX2X1_1 MUX2X1_1/A MUX2X1_1/B MUX2X1_1/S gnd MUX2X1_1/Y vdd MUX2X1
XCLKBUF1_2 CLKBUF1_8/A gnd CLKBUF1_2/Y vdd CLKBUF1
XBUFX4_162 wb_sel_i[2] gnd BUFX4_162/Y vdd BUFX4
XBUFX4_151 BUFX4_152/A gnd BUFX4_151/Y vdd BUFX4
XBUFX4_140 INVX8_7/Y gnd DFFSR_53/R vdd BUFX4
XNOR2X1_211 NOR2X1_243/B INVX8_14/Y gnd NOR2X1_211/Y vdd NOR2X1
XBUFX4_184 BUFX4_185/A gnd BUFX4_184/Y vdd BUFX4
XNOR2X1_233 DFFSR_209/Q BUFX4_35/Y gnd NOR2X1_233/Y vdd NOR2X1
XNOR2X1_222 NOR2X1_238/B OR2X2_12/A gnd NOR2X1_222/Y vdd NOR2X1
XBUFX4_195 BUFX4_194/A gnd BUFX4_195/Y vdd BUFX4
XNOR2X1_200 miso_pad_i INVX1_121/Y gnd NOR2X1_200/Y vdd NOR2X1
XBUFX4_173 BUFX4_172/A gnd BUFX4_173/Y vdd BUFX4
XOAI21X1_717 NOR2X1_320/Y OAI21X1_716/Y OAI21X1_717/C gnd DFFSR_121/D vdd OAI21X1
XOAI21X1_728 NOR2X1_322/Y OAI21X1_728/B NAND2X1_322/Y gnd DFFSR_118/D vdd OAI21X1
XNOR2X1_244 INVX2_55/A BUFX4_36/Y gnd NOR2X1_244/Y vdd NOR2X1
XNOR2X1_277 INVX2_88/A BUFX4_115/Y gnd NOR2X1_277/Y vdd NOR2X1
XNOR2X1_288 INVX1_47/A BUFX4_115/Y gnd NOR2X1_288/Y vdd NOR2X1
XOAI21X1_739 BUFX4_168/Y OAI21X1_738/Y BUFX4_38/Y gnd OAI21X1_740/B vdd OAI21X1
XNOR2X1_255 INVX2_63/A BUFX4_38/Y gnd NOR2X1_255/Y vdd NOR2X1
XNOR2X1_299 INVX8_22/Y OR2X2_18/A gnd INVX1_143/A vdd NOR2X1
XNOR2X1_266 BUFX4_229/Y OR2X2_14/A gnd NOR2X1_266/Y vdd NOR2X1
XOAI21X1_706 OAI21X1_706/A BUFX4_210/Y OAI21X1_706/C gnd DFFSR_125/D vdd OAI21X1
XINVX8_4 INVX8_4/A gnd INVX8_4/Y vdd INVX8
XBUFX4_24 INVX8_1/Y gnd BUFX4_24/Y vdd BUFX4
XBUFX4_79 wb_sel_i[0] gnd BUFX4_79/Y vdd BUFX4
XBUFX4_13 BUFX4_19/A gnd AND2X2_2/B vdd BUFX4
XBUFX4_68 wb_sel_i[3] gnd MUX2X1_7/S vdd BUFX4
XBUFX4_46 BUFX4_45/A gnd BUFX4_46/Y vdd BUFX4
XBUFX4_35 BUFX4_36/A gnd BUFX4_35/Y vdd BUFX4
XBUFX4_57 BUFX4_61/A gnd BUFX4_57/Y vdd BUFX4
XFILL_30_2_0 gnd vdd FILL
XOR2X2_9 OR2X2_9/A OR2X2_9/B gnd OR2X2_9/Y vdd OR2X2
XOR2X2_16 OR2X2_16/A INVX4_9/Y gnd OR2X2_16/Y vdd OR2X2
XINVX2_162 DFFSR_233/Q gnd INVX2_162/Y vdd INVX2
XINVX2_151 INVX2_151/A gnd INVX2_151/Y vdd INVX2
XINVX2_140 INVX1_48/A gnd MUX2X1_3/A vdd INVX2
XINVX8_16 BUFX4_50/Y gnd INVX8_16/Y vdd INVX8
XOAI21X1_547 OAI21X1_547/A OAI21X1_547/B OAI21X1_543/Y gnd DFFSR_182/D vdd OAI21X1
XOAI21X1_525 INVX2_59/Y BUFX4_85/Y NAND2X1_239/Y gnd OAI21X1_525/Y vdd OAI21X1
XFILL_21_2_0 gnd vdd FILL
XOAI21X1_536 BUFX4_169/Y OAI21X1_535/Y BUFX4_37/Y gnd OAI21X1_537/B vdd OAI21X1
XOAI21X1_558 AND2X2_28/Y INVX2_64/Y BUFX4_119/Y gnd OAI21X1_558/Y vdd OAI21X1
XOAI21X1_569 OAI21X1_569/A OAI21X1_569/B NAND2X1_260/Y gnd DFFSR_175/D vdd OAI21X1
XOAI21X1_503 NOR2X1_257/Y INVX2_86/Y BUFX4_166/Y gnd OAI21X1_503/Y vdd OAI21X1
XOAI21X1_514 AND2X2_24/Y MUX2X1_4/A BUFX4_166/Y gnd AOI21X1_180/C vdd OAI21X1
XFILL_29_3_0 gnd vdd FILL
XFILL_4_3_0 gnd vdd FILL
XFILL_12_2_0 gnd vdd FILL
XNAND3X1_181 INVX2_49/Y NAND3X1_180/Y NAND2X1_143/B gnd AND2X2_20/B vdd NAND3X1
XNAND3X1_170 INVX2_43/A OR2X2_8/A OR2X2_8/B gnd INVX1_103/A vdd NAND3X1
XNAND3X1_192 AND2X2_20/Y AOI21X1_43/Y AOI21X1_45/B gnd NAND3X1_193/C vdd NAND3X1
XOAI21X1_311 INVX2_73/A BUFX4_176/Y AOI21X1_97/Y gnd NAND3X1_207/B vdd OAI21X1
XOAI21X1_377 INVX2_148/Y BUFX4_165/Y NAND2X1_226/Y gnd OAI21X1_377/Y vdd OAI21X1
XOAI21X1_366 BUFX4_59/Y NAND2X1_218/Y OAI21X1_366/C gnd OAI21X1_366/Y vdd OAI21X1
XOAI21X1_333 INVX2_81/Y BUFX4_70/Y OAI21X1_333/C gnd OAI21X1_333/Y vdd OAI21X1
XOAI21X1_399 BUFX4_55/Y OAI21X1_399/B BUFX4_240/Y gnd OAI21X1_399/Y vdd OAI21X1
XOAI21X1_344 BUFX4_55/Y OAI21X1_343/Y BUFX4_240/Y gnd OAI21X1_345/B vdd OAI21X1
XOAI21X1_322 AND2X2_22/Y INVX2_65/Y BUFX4_53/Y gnd OAI21X1_322/Y vdd OAI21X1
XOAI21X1_355 OAI21X1_355/A OAI21X1_354/Y OAI21X1_355/C gnd DFFSR_236/D vdd OAI21X1
XOAI21X1_300 INVX2_83/A BUFX4_177/Y AOI21X1_74/Y gnd OAI21X1_300/Y vdd OAI21X1
XOAI21X1_388 OAI21X1_388/A OAI21X1_388/B OAI21X1_384/Y gnd DFFSR_225/D vdd OAI21X1
XDFFSR_190 INVX2_72/A CLKBUF1_34/Y DFFSR_167/R vdd DFFSR_190/D gnd vdd DFFSR
XFILL_35_1_0 gnd vdd FILL
XNAND3X1_1 wb_stb_i wb_cyc_i wb_we_i gnd NOR2X1_1/B vdd NAND3X1
XFILL_27_6_1 gnd vdd FILL
XFILL_26_1_0 gnd vdd FILL
XFILL_2_6_1 gnd vdd FILL
XFILL_1_1_0 gnd vdd FILL
XOAI21X1_130 BUFX4_95/Y BUFX4_102/Y DFFSR_4/Q gnd BUFX2_6/A vdd OAI21X1
XFILL_10_5_1 gnd vdd FILL
XAOI22X1_6 INVX2_78/A AOI22X1_1/B INVX8_6/Y INVX2_77/A gnd AOI22X1_6/Y vdd AOI22X1
XOAI21X1_196 AND2X2_11/Y NOR2X1_63/Y BUFX4_245/Y gnd OAI21X1_197/C vdd OAI21X1
XOAI21X1_141 BUFX4_95/Y BUFX4_102/Y INVX2_7/A gnd BUFX2_17/A vdd OAI21X1
XOAI21X1_185 INVX1_83/Y NOR2X1_54/Y INVX8_9/A gnd OAI21X1_186/C vdd OAI21X1
XOAI21X1_152 BUFX4_94/Y BUFX4_97/Y INVX1_2/A gnd BUFX2_28/A vdd OAI21X1
XOAI21X1_174 XNOR2X1_2/Y BUFX4_2/Y NAND2X1_97/Y gnd DFFSR_109/D vdd OAI21X1
XOAI21X1_163 XOR2X1_1/A XOR2X1_1/B INVX1_70/A gnd AND2X2_6/B vdd OAI21X1
XNAND2X1_16 NAND2X1_9/B wb_dat_i[23] gnd OAI21X1_31/C vdd NAND2X1
XNAND2X1_27 BUFX4_83/Y wb_dat_i[2] gnd NAND2X1_27/Y vdd NAND2X1
XNAND2X1_38 NAND3X1_71/Y NAND3X1_72/Y gnd AOI21X1_2/C vdd NAND2X1
XNAND2X1_49 AOI21X1_9/Y NOR2X1_12/Y gnd DFFSR_73/D vdd NAND2X1
XNAND2X1_180 INVX2_88/Y BUFX4_175/Y gnd AOI22X1_52/A vdd NAND2X1
XNAND2X1_191 AOI22X1_62/Y AOI22X1_63/Y gnd NAND2X1_191/Y vdd NAND2X1
XFILL_9_2_0 gnd vdd FILL
XFILL_18_6_1 gnd vdd FILL
XFILL_17_1_0 gnd vdd FILL
XAOI22X1_36 AOI22X1_36/A AOI21X1_32/Y AOI22X1_36/C INVX1_115/A gnd BUFX4_172/A vdd
+ AOI22X1
XAOI22X1_14 BUFX4_25/Y INVX1_15/A INVX2_52/A INVX8_6/Y gnd AOI22X1_14/Y vdd AOI22X1
XAOI22X1_47 AOI22X1_47/A AOI21X1_69/Y AOI22X1_47/C AOI22X1_47/D gnd AOI22X1_47/Y vdd
+ AOI22X1
XAOI21X1_209 AOI21X1_209/A AOI21X1_209/B NOR2X1_279/Y gnd DFFSR_167/D vdd AOI21X1
XAOI22X1_25 INVX2_82/A BUFX4_124/Y INVX8_5/Y INVX2_83/A gnd NAND3X1_98/B vdd AOI22X1
XAOI22X1_69 INVX2_64/A INVX4_9/A INVX4_7/A INVX2_66/A gnd AOI22X1_69/Y vdd AOI22X1
XAOI22X1_58 DFFSR_243/Q INVX8_14/A INVX8_22/A AND2X2_17/B gnd AOI22X1_58/Y vdd AOI22X1
XOAI22X1_9 OAI22X1_9/A INVX1_34/Y INVX8_2/A INVX2_19/Y gnd AOI21X1_4/C vdd OAI22X1
XAOI21X1_91 INVX2_132/Y BUFX4_156/Y AOI21X1_69/C gnd AOI22X1_56/D vdd AOI21X1
XAOI21X1_80 INVX2_90/Y BUFX4_175/Y INVX1_118/A gnd AOI21X1_80/Y vdd AOI21X1
XFILL_33_4_1 gnd vdd FILL
XINVX2_18 INVX2_18/A gnd INVX2_18/Y vdd INVX2
XINVX2_29 INVX2_29/A gnd INVX2_29/Y vdd INVX2
XFILL_24_4_1 gnd vdd FILL
XFILL_6_0_0 gnd vdd FILL
XFILL_7_5_1 gnd vdd FILL
XXOR2X1_1 XOR2X1_1/A XOR2X1_1/B gnd XOR2X1_1/Y vdd XOR2X1
XFILL_15_4_1 gnd vdd FILL
XMUX2X1_2 MUX2X1_2/A MUX2X1_2/B MUX2X1_1/S gnd MUX2X1_2/Y vdd MUX2X1
XCLKBUF1_3 CLKBUF1_3/A gnd DFFSR_5/CLK vdd CLKBUF1
XBUFX4_130 INVX8_24/Y gnd BUFX4_130/Y vdd BUFX4
XBUFX4_163 wb_sel_i[2] gnd BUFX4_163/Y vdd BUFX4
XFILL_31_1 gnd vdd FILL
XBUFX4_152 BUFX4_152/A gnd BUFX4_152/Y vdd BUFX4
XBUFX4_185 BUFX4_185/A gnd BUFX4_185/Y vdd BUFX4
XNOR2X1_245 BUFX4_150/Y NOR2X1_245/B gnd AND2X2_26/A vdd NOR2X1
XNOR2X1_234 BUFX4_96/Y INVX1_132/Y gnd BUFX4_211/A vdd NOR2X1
XBUFX4_141 INVX8_7/Y gnd DFFSR_58/R vdd BUFX4
XBUFX4_174 BUFX4_172/A gnd BUFX4_174/Y vdd BUFX4
XNOR2X1_212 NOR2X1_245/B INVX8_14/Y gnd NOR2X1_212/Y vdd NOR2X1
XNOR2X1_267 INVX2_151/A BUFX4_116/Y gnd NOR2X1_267/Y vdd NOR2X1
XBUFX4_196 BUFX4_194/A gnd AND2X2_16/B vdd BUFX4
XNOR2X1_223 NOR2X1_239/B OR2X2_12/A gnd NOR2X1_223/Y vdd NOR2X1
XNOR2X1_256 INVX4_8/Y OR2X2_14/A gnd NOR2X1_256/Y vdd NOR2X1
XNOR2X1_201 BUFX4_99/Y INVX4_6/Y gnd BUFX4_152/A vdd NOR2X1
XOAI21X1_729 INVX1_99/Y BUFX4_80/Y NAND2X1_245/Y gnd OAI21X1_729/Y vdd OAI21X1
XNOR2X1_289 INVX1_41/A BUFX4_115/Y gnd NOR2X1_289/Y vdd NOR2X1
XOAI21X1_718 INVX2_94/Y BUFX4_85/Y NAND2X1_242/Y gnd OAI21X1_718/Y vdd OAI21X1
XNOR2X1_278 INVX8_19/A NOR2X1_262/B gnd NOR2X1_278/Y vdd NOR2X1
XOAI21X1_707 INVX2_96/Y BUFX4_5/Y NAND2X1_238/Y gnd NAND2X1_313/B vdd OAI21X1
XINVX8_5 INVX8_5/A gnd INVX8_5/Y vdd INVX8
XBUFX4_25 INVX8_1/Y gnd BUFX4_25/Y vdd BUFX4
XBUFX4_14 BUFX4_19/A gnd BUFX4_14/Y vdd BUFX4
XBUFX4_36 BUFX4_36/A gnd BUFX4_36/Y vdd BUFX4
XBUFX4_58 BUFX4_61/A gnd BUFX4_58/Y vdd BUFX4
XBUFX4_47 BUFX4_47/A gnd BUFX4_47/Y vdd BUFX4
XBUFX4_69 wb_sel_i[3] gnd MUX2X1_8/S vdd BUFX4
XFILL_30_2_1 gnd vdd FILL
XINVX2_163 DFFSR_169/Q gnd INVX2_163/Y vdd INVX2
XOR2X2_17 OR2X2_17/A OR2X2_17/B gnd OR2X2_17/Y vdd OR2X2
XINVX2_130 INVX2_130/A gnd INVX2_130/Y vdd INVX2
XINVX2_141 INVX2_141/A gnd MUX2X1_3/B vdd INVX2
XINVX2_152 DFFSR_209/Q gnd INVX2_152/Y vdd INVX2
XINVX8_17 INVX8_17/A gnd OR2X2_12/A vdd INVX8
XOAI21X1_548 BUFX4_211/Y BUFX4_32/Y INVX2_146/A gnd OAI21X1_552/C vdd OAI21X1
XOAI21X1_526 BUFX4_170/Y OAI21X1_525/Y BUFX4_37/Y gnd OAI21X1_527/B vdd OAI21X1
XFILL_21_2_1 gnd vdd FILL
XOAI21X1_537 OAI21X1_537/A OAI21X1_537/B OAI21X1_533/Y gnd DFFSR_184/D vdd OAI21X1
XOAI21X1_559 INVX2_64/Y BUFX4_72/Y OAI21X1_323/C gnd OAI21X1_560/B vdd OAI21X1
XOAI21X1_504 INVX2_86/Y BUFX4_11/Y OAI21X1_699/C gnd OAI21X1_505/B vdd OAI21X1
XOAI21X1_515 MUX2X1_4/A BUFX4_6/Y OAI21X1_515/C gnd OAI21X1_516/B vdd OAI21X1
XFILL_29_3_1 gnd vdd FILL
XFILL_4_3_1 gnd vdd FILL
XFILL_12_2_1 gnd vdd FILL
XNAND3X1_160 INVX8_10/Y OAI21X1_257/Y NAND3X1_160/C gnd NAND3X1_162/B vdd NAND3X1
XNAND3X1_171 INVX2_48/Y BUFX4_111/Y INVX1_103/Y gnd NAND2X1_129/B vdd NAND3X1
XNAND3X1_182 AOI21X1_43/A NAND2X1_144/B AOI21X1_37/Y gnd NAND3X1_182/Y vdd NAND3X1
XNAND3X1_193 BUFX4_248/Y NAND3X1_185/C NAND3X1_193/C gnd AND2X2_21/A vdd NAND3X1
XOAI21X1_312 INVX2_55/A BUFX4_176/Y AOI21X1_100/Y gnd NAND3X1_208/A vdd OAI21X1
XOAI21X1_323 INVX2_65/Y BUFX4_73/Y OAI21X1_323/C gnd OAI21X1_323/Y vdd OAI21X1
XOAI21X1_301 DFFSR_172/Q BUFX4_158/Y AOI21X1_83/Y gnd OAI21X1_301/Y vdd OAI21X1
XDFFSR_180 DFFSR_180/Q CLKBUF1_54/Y DFFSR_165/R vdd DFFSR_180/D gnd vdd DFFSR
XOAI21X1_367 INVX2_89/Y NAND2X1_9/B NAND2X1_219/Y gnd OAI21X1_367/Y vdd OAI21X1
XOAI21X1_378 BUFX4_52/Y OAI21X1_377/Y BUFX4_241/Y gnd OAI21X1_378/Y vdd OAI21X1
XOAI21X1_356 BUFX4_220/Y BUFX4_230/Y INVX2_52/A gnd OAI21X1_356/Y vdd OAI21X1
XOAI21X1_334 BUFX4_55/Y OAI21X1_333/Y BUFX4_240/Y gnd OAI21X1_335/B vdd OAI21X1
XOAI21X1_345 OAI21X1_345/A OAI21X1_345/B OAI21X1_341/Y gnd DFFSR_238/D vdd OAI21X1
XDFFSR_191 INVX1_53/A CLKBUF1_32/Y DFFSR_167/R vdd DFFSR_191/D gnd vdd DFFSR
XOAI21X1_389 BUFX4_222/Y BUFX4_233/Y INVX1_55/A gnd OAI21X1_389/Y vdd OAI21X1
XNAND2X1_340 BUFX4_206/Y OAI21X1_787/Y gnd NAND2X1_340/Y vdd NAND2X1
XFILL_35_1_1 gnd vdd FILL
XNAND3X1_2 wb_adr_i[4] wb_adr_i[3] INVX4_1/Y gnd BUFX4_78/A vdd NAND3X1
XFILL_26_1_1 gnd vdd FILL
XFILL_1_1_1 gnd vdd FILL
XOAI21X1_131 BUFX4_93/Y BUFX4_103/Y DFFSR_5/Q gnd BUFX2_7/A vdd OAI21X1
XOAI21X1_120 INVX2_36/Y BUFX4_84/Y OAI21X1_59/C gnd NAND3X1_64/B vdd OAI21X1
XAOI22X1_7 AOI22X1_7/A AOI22X1_7/B INVX8_5/Y DFFSR_199/Q gnd AOI22X1_7/Y vdd AOI22X1
XOAI21X1_153 BUFX4_91/Y BUFX4_97/Y INVX1_3/A gnd BUFX2_29/A vdd OAI21X1
XOAI21X1_142 BUFX4_94/Y NOR2X1_1/A INVX2_8/A gnd BUFX2_18/A vdd OAI21X1
XOAI21X1_164 BUFX4_1/Y AND2X2_6/Y NAND2X1_90/Y gnd DFFSR_102/D vdd OAI21X1
XOAI21X1_197 BUFX4_248/Y NAND2X1_107/Y OAI21X1_197/C gnd BUFX4_239/A vdd OAI21X1
XOAI21X1_186 INVX8_9/A INVX2_45/Y OAI21X1_186/C gnd INVX1_84/A vdd OAI21X1
XOAI21X1_175 AND2X2_8/Y AOI21X1_23/Y NOR2X1_46/B gnd OAI21X1_176/C vdd OAI21X1
XFILL_9_2_1 gnd vdd FILL
XNAND2X1_39 AOI21X1_2/Y NOR2X1_5/Y gnd DFFSR_66/D vdd NAND2X1
XNAND2X1_28 BUFX4_85/Y wb_dat_i[3] gnd NAND2X1_28/Y vdd NAND2X1
XNAND2X1_170 INVX1_17/A INVX1_80/Y gnd NAND2X1_170/Y vdd NAND2X1
XNAND2X1_17 wb_dat_i[8] BUFX4_5/Y gnd OAI21X1_33/C vdd NAND2X1
XNAND2X1_181 INVX2_91/Y BUFX4_155/Y gnd AOI22X1_52/D vdd NAND2X1
XNAND2X1_192 AOI22X1_64/Y AOI22X1_65/Y gnd NAND2X1_192/Y vdd NAND2X1
XFILL_17_1_1 gnd vdd FILL
XAOI22X1_48 AOI22X1_48/A AOI21X1_71/Y AOI21X1_72/Y AOI22X1_48/D gnd AOI22X1_48/Y vdd
+ AOI22X1
XAOI22X1_15 BUFX4_25/Y INVX1_16/A INVX2_130/A INVX8_5/Y gnd AOI22X1_15/Y vdd AOI22X1
XAOI22X1_37 AOI22X1_37/A AOI22X1_37/B AOI22X1_37/C INVX1_117/Y gnd AOI22X1_37/Y vdd
+ AOI22X1
XAOI22X1_26 BUFX4_22/Y INVX1_5/A INVX2_81/A INVX8_6/Y gnd NAND3X1_98/C vdd AOI22X1
XAOI22X1_59 INVX1_62/A INVX8_17/A INVX4_7/A INVX2_127/A gnd AOI22X1_59/Y vdd AOI22X1
XAOI21X1_70 INVX2_107/Y BUFX4_172/Y INVX1_117/A gnd AOI22X1_47/C vdd AOI21X1
XAOI21X1_92 INVX2_131/Y BUFX4_174/Y INVX1_118/A gnd AOI21X1_92/Y vdd AOI21X1
XAOI21X1_81 INVX2_99/Y BUFX4_153/Y AOI21X1_69/C gnd AOI22X1_53/B vdd AOI21X1
XINVX2_19 INVX4_3/A gnd INVX2_19/Y vdd INVX2
XXOR2X1_2 XOR2X1_2/A XOR2X1_2/B gnd XOR2X1_2/Y vdd XOR2X1
XFILL_6_0_1 gnd vdd FILL
XMUX2X1_3 MUX2X1_3/A MUX2X1_3/B MUX2X1_1/S gnd MUX2X1_3/Y vdd MUX2X1
XCLKBUF1_4 CLKBUF1_4/A gnd CLKBUF1_4/Y vdd CLKBUF1
XBUFX4_120 INVX8_20/Y gnd BUFX4_120/Y vdd BUFX4
XBUFX4_197 BUFX4_194/A gnd BUFX4_197/Y vdd BUFX4
XBUFX4_164 wb_sel_i[2] gnd BUFX4_164/Y vdd BUFX4
XNOR2X1_213 INVX2_89/A BUFX4_241/Y gnd NOR2X1_213/Y vdd NOR2X1
XFILL_24_1 gnd vdd FILL
XBUFX4_142 INVX8_7/Y gnd DFFSR_9/R vdd BUFX4
XNOR2X1_246 INVX2_160/A BUFX4_39/Y gnd NOR2X1_246/Y vdd NOR2X1
XNOR2X1_279 AOI22X1_7/A BUFX4_115/Y gnd NOR2X1_279/Y vdd NOR2X1
XBUFX4_186 BUFX4_185/A gnd AND2X2_15/B vdd BUFX4
XBUFX4_131 INVX8_24/Y gnd DFFSR_167/R vdd BUFX4
XNOR2X1_268 BUFX4_229/Y NOR2X1_257/B gnd AND2X2_30/A vdd NOR2X1
XNOR2X1_235 BUFX4_96/Y INVX8_18/Y gnd BUFX4_32/A vdd NOR2X1
XNOR2X1_202 INVX1_122/Y INVX2_164/Y gnd AND2X2_22/A vdd NOR2X1
XNOR2X1_257 INVX4_8/Y NOR2X1_257/B gnd NOR2X1_257/Y vdd NOR2X1
XNOR2X1_224 NOR2X1_224/A OR2X2_12/A gnd NOR2X1_224/Y vdd NOR2X1
XBUFX4_153 BUFX4_154/A gnd BUFX4_153/Y vdd BUFX4
XBUFX4_175 BUFX4_172/A gnd BUFX4_175/Y vdd BUFX4
XOAI21X1_719 INVX1_150/A OR2X2_18/B INVX2_94/Y gnd OAI21X1_720/C vdd OAI21X1
XOAI21X1_708 OR2X2_19/A OR2X2_18/B INVX2_96/Y gnd OAI21X1_709/C vdd OAI21X1
XINVX8_6 INVX8_6/A gnd INVX8_6/Y vdd INVX8
XBUFX4_26 INVX8_1/Y gnd BUFX4_26/Y vdd BUFX4
XBUFX4_15 BUFX4_19/A gnd BUFX4_15/Y vdd BUFX4
XBUFX4_48 BUFX4_47/A gnd BUFX4_48/Y vdd BUFX4
XBUFX4_37 BUFX4_36/A gnd BUFX4_37/Y vdd BUFX4
XBUFX4_59 BUFX4_61/A gnd BUFX4_59/Y vdd BUFX4
XINVX2_131 DFFSR_139/Q gnd INVX2_131/Y vdd INVX2
XINVX2_120 AOI22X1_8/C gnd INVX2_120/Y vdd INVX2
XOR2X2_18 OR2X2_18/A OR2X2_18/B gnd OR2X2_18/Y vdd OR2X2
XINVX2_153 INVX1_59/A gnd INVX2_153/Y vdd INVX2
XINVX2_164 INVX2_164/A gnd INVX2_164/Y vdd INVX2
XINVX2_142 DFFSR_189/Q gnd MUX2X1_4/A vdd INVX2
XINVX8_18 INVX8_18/A gnd INVX8_18/Y vdd INVX8
XOAI21X1_505 BUFX4_167/Y OAI21X1_505/B BUFX4_39/Y gnd OAI21X1_506/B vdd OAI21X1
XOAI21X1_549 NOR2X1_264/Y INVX2_146/Y BUFX4_171/Y gnd AOI21X1_187/C vdd OAI21X1
XOAI21X1_527 AOI21X1_182/Y OAI21X1_527/B OAI21X1_523/Y gnd DFFSR_186/D vdd OAI21X1
XOAI21X1_538 INVX8_21/A BUFX4_28/Y INVX1_33/A gnd OAI21X1_542/C vdd OAI21X1
XOAI21X1_516 BUFX4_166/Y OAI21X1_516/B BUFX4_39/Y gnd OAI21X1_517/B vdd OAI21X1
XAOI21X1_190 INVX2_151/Y NAND2X1_258/Y BUFX4_29/Y gnd AOI21X1_190/Y vdd AOI21X1
XFILL_31_5_0 gnd vdd FILL
XNAND3X1_150 INVX4_4/Y NAND3X1_148/Y NAND3X1_149/Y gnd NAND3X1_150/Y vdd NAND3X1
XNAND3X1_183 INVX1_116/A INVX1_105/A NAND3X1_182/Y gnd INVX1_115/A vdd NAND3X1
XNAND3X1_172 INVX2_46/Y AOI21X1_33/A AOI21X1_33/B gnd AOI21X1_34/B vdd NAND3X1
XNAND3X1_194 INVX1_106/Y NAND2X1_149/Y NAND3X1_191/Y gnd AOI21X1_71/C vdd NAND3X1
XNAND3X1_161 BUFX4_237/Y NAND3X1_161/B OAI21X1_260/Y gnd NAND3X1_161/Y vdd NAND3X1
XOAI21X1_313 INVX1_42/A BUFX4_178/Y AOI21X1_101/Y gnd OAI21X1_313/Y vdd OAI21X1
XFILL_22_5_0 gnd vdd FILL
XOAI21X1_346 BUFX4_224/Y BUFX4_231/Y INVX2_141/A gnd OAI21X1_350/C vdd OAI21X1
XOAI21X1_335 OAI21X1_335/A OAI21X1_335/B OAI21X1_331/Y gnd DFFSR_240/D vdd OAI21X1
XOAI21X1_324 BUFX4_53/Y OAI21X1_323/Y BUFX4_242/Y gnd OAI21X1_324/Y vdd OAI21X1
XOAI21X1_302 DFFSR_204/Q BUFX4_177/Y AOI21X1_84/Y gnd OAI21X1_302/Y vdd OAI21X1
XDFFSR_170 INVX2_54/A CLKBUF1_4/Y DFFSR_165/R vdd DFFSR_170/D gnd vdd DFFSR
XOAI21X1_379 AOI21X1_120/Y OAI21X1_378/Y OAI21X1_379/C gnd DFFSR_229/D vdd OAI21X1
XDFFSR_181 INVX2_146/A CLKBUF1_19/Y DFFSR_137/R vdd DFFSR_181/D gnd vdd DFFSR
XOAI21X1_357 NOR2X1_211/Y INVX2_52/Y BUFX4_52/Y gnd AOI21X1_111/C vdd OAI21X1
XOAI21X1_368 BUFX4_59/Y NAND2X1_221/Y OAI21X1_368/C gnd AOI21X1_118/B vdd OAI21X1
XDFFSR_192 INVX2_86/A CLKBUF1_28/Y DFFSR_167/R vdd DFFSR_192/D gnd vdd DFFSR
XNAND2X1_330 BUFX4_161/Y wb_dat_i[23] gnd NAND2X1_330/Y vdd NAND2X1
XNAND2X1_341 INVX8_23/A INVX1_164/A gnd OAI21X1_789/B vdd NAND2X1
XFILL_5_6_0 gnd vdd FILL
XFILL_13_5_0 gnd vdd FILL
XNAND3X1_3 BUFX4_14/Y OAI21X1_1/Y BUFX4_22/Y gnd OAI21X1_2/C vdd NAND3X1
XOAI21X1_198 INVX1_86/Y INVX2_42/A OR2X2_7/B gnd NAND2X1_108/A vdd OAI21X1
XOAI21X1_143 BUFX4_92/Y INVX4_5/A INVX1_9/A gnd BUFX2_19/A vdd OAI21X1
XOAI21X1_132 BUFX4_93/Y BUFX4_103/Y DFFSR_6/Q gnd BUFX2_8/A vdd OAI21X1
XOAI21X1_187 OR2X2_8/A OR2X2_8/B INVX2_43/A gnd OAI21X1_187/Y vdd OAI21X1
XOAI21X1_110 INVX2_31/Y BUFX4_79/Y NAND2X1_25/Y gnd NAND3X1_59/B vdd OAI21X1
XOAI21X1_121 AND2X2_3/Y INVX2_36/Y NAND3X1_64/Y gnd DFFSR_52/D vdd OAI21X1
XAOI22X1_8 BUFX4_25/Y DFFSR_20/Q AOI22X1_8/C INVX8_6/Y gnd AOI22X1_8/Y vdd AOI22X1
XOAI21X1_154 BUFX4_94/Y BUFX4_97/Y INVX1_4/A gnd BUFX2_30/A vdd OAI21X1
XOAI21X1_176 INVX1_68/Y NOR2X1_46/B OAI21X1_176/C gnd DFFSR_110/D vdd OAI21X1
XOAI21X1_165 BUFX4_3/Y AOI21X1_20/Y NAND2X1_91/Y gnd DFFSR_103/D vdd OAI21X1
XNAND2X1_29 BUFX4_79/Y wb_dat_i[4] gnd OAI21X1_86/C vdd NAND2X1
XNAND2X1_171 INVX2_105/Y BUFX4_172/Y gnd AOI22X1_47/A vdd NAND2X1
XNAND2X1_193 INVX2_78/Y BUFX4_178/Y gnd AOI22X1_66/B vdd NAND2X1
XNAND2X1_182 AOI22X1_51/Y AOI22X1_52/Y gnd AOI22X1_54/B vdd NAND2X1
XNAND2X1_160 AOI22X1_39/Y AOI22X1_40/Y gnd AOI22X1_41/D vdd NAND2X1
XNAND2X1_18 BUFX4_7/Y wb_dat_i[9] gnd OAI21X1_65/C vdd NAND2X1
XAOI22X1_38 AOI21X1_55/Y AOI22X1_38/B AOI22X1_38/C INVX1_118/Y gnd AOI22X1_38/Y vdd
+ AOI22X1
XAOI22X1_16 INVX2_129/A AOI22X1_7/B INVX8_6/Y INVX2_128/A gnd AOI22X1_16/Y vdd AOI22X1
XAOI22X1_27 INVX8_6/Y INVX2_150/A DFFSR_209/Q INVX8_5/Y gnd NAND3X1_99/C vdd AOI22X1
XAOI22X1_49 AOI21X1_76/Y AOI22X1_49/B AOI22X1_49/C AOI22X1_49/D gnd AOI22X1_49/Y vdd
+ AOI22X1
XFILL_27_4_0 gnd vdd FILL
XFILL_2_4_0 gnd vdd FILL
XAOI21X1_71 INVX2_102/Y BUFX4_154/Y AOI21X1_71/C gnd AOI21X1_71/Y vdd AOI21X1
XAOI21X1_60 INVX2_158/Y BUFX4_157/Y AOI21X1_69/C gnd AOI21X1_60/Y vdd AOI21X1
XAOI21X1_93 INVX2_135/Y BUFX4_178/Y INVX1_117/A gnd AOI21X1_93/Y vdd AOI21X1
XFILL_10_3_0 gnd vdd FILL
XAOI21X1_82 INVX2_96/Y BUFX4_173/Y INVX1_117/A gnd AOI21X1_82/Y vdd AOI21X1
XFILL_18_4_0 gnd vdd FILL
XXOR2X1_3 XOR2X1_3/A XOR2X1_3/B gnd OR2X2_9/B vdd XOR2X1
XMUX2X1_4 MUX2X1_4/A MUX2X1_4/B MUX2X1_1/S gnd MUX2X1_4/Y vdd MUX2X1
XCLKBUF1_5 CLKBUF1_5/A gnd CLKBUF1_5/Y vdd CLKBUF1
XBUFX4_110 DFFSR_42/Q gnd INVX8_13/A vdd BUFX4
XBUFX4_132 INVX8_24/Y gnd DFFSR_165/R vdd BUFX4
XBUFX4_121 INVX8_20/Y gnd BUFX4_121/Y vdd BUFX4
XBUFX4_154 BUFX4_154/A gnd BUFX4_154/Y vdd BUFX4
XBUFX4_143 INVX8_7/Y gnd DFFSR_25/R vdd BUFX4
XFILL_33_2_0 gnd vdd FILL
XBUFX4_165 wb_sel_i[2] gnd BUFX4_165/Y vdd BUFX4
XFILL_24_2 gnd vdd FILL
XBUFX4_176 BUFX4_172/A gnd BUFX4_176/Y vdd BUFX4
XNOR2X1_225 NOR2X1_243/B OR2X2_12/A gnd NOR2X1_225/Y vdd NOR2X1
XNOR2X1_214 AOI22X1_8/C BUFX4_244/Y gnd NOR2X1_214/Y vdd NOR2X1
XFILL_17_1 gnd vdd FILL
XNOR2X1_247 INVX2_91/A BUFX4_39/Y gnd NOR2X1_247/Y vdd NOR2X1
XNOR2X1_269 INVX2_82/A BUFX4_116/Y gnd NOR2X1_269/Y vdd NOR2X1
XBUFX4_198 BUFX4_194/A gnd BUFX4_198/Y vdd BUFX4
XNOR2X1_258 INVX1_53/A BUFX4_38/Y gnd NOR2X1_258/Y vdd NOR2X1
XNOR2X1_236 INVX4_7/Y NOR2X1_257/B gnd NOR2X1_236/Y vdd NOR2X1
XBUFX4_187 BUFX4_185/A gnd BUFX4_187/Y vdd BUFX4
XNOR2X1_203 INVX1_125/A INVX2_164/Y gnd INVX1_123/A vdd NOR2X1
XOAI21X1_709 BUFX4_62/Y OR2X2_19/Y OAI21X1_709/C gnd OAI21X1_710/A vdd OAI21X1
XFILL_24_2_0 gnd vdd FILL
XINVX8_7 wb_rst_i gnd INVX8_7/Y vdd INVX8
XBUFX4_16 BUFX4_19/A gnd BUFX4_16/Y vdd BUFX4
XBUFX4_27 INVX8_1/Y gnd BUFX4_27/Y vdd BUFX4
XBUFX4_49 BUFX4_47/A gnd BUFX4_49/Y vdd BUFX4
XBUFX4_38 BUFX4_36/A gnd BUFX4_38/Y vdd BUFX4
XFILL_7_3_0 gnd vdd FILL
XFILL_15_2_0 gnd vdd FILL
XINVX2_132 INVX1_44/A gnd INVX2_132/Y vdd INVX2
XINVX2_121 AOI22X1_7/A gnd INVX2_121/Y vdd INVX2
XINVX2_110 INVX2_110/A gnd INVX2_110/Y vdd INVX2
XOR2X2_19 OR2X2_19/A OR2X2_18/B gnd OR2X2_19/Y vdd OR2X2
XINVX2_143 DFFSR_205/Q gnd MUX2X1_4/B vdd INVX2
XINVX2_165 INVX2_165/A gnd INVX2_165/Y vdd INVX2
XINVX2_154 INVX1_57/A gnd INVX2_154/Y vdd INVX2
XOAI21X1_528 INVX8_21/A BUFX4_33/Y INVX1_39/A gnd OAI21X1_528/Y vdd OAI21X1
XOAI21X1_539 NOR2X1_262/Y INVX2_116/Y BUFX4_169/Y gnd AOI21X1_185/C vdd OAI21X1
XINVX8_19 INVX8_19/A gnd INVX8_19/Y vdd INVX8
XOAI21X1_506 OAI21X1_506/A OAI21X1_506/B OAI21X1_502/Y gnd DFFSR_192/D vdd OAI21X1
XOAI21X1_517 OAI21X1_517/A OAI21X1_517/B OAI21X1_513/Y gnd DFFSR_189/D vdd OAI21X1
XAOI21X1_191 BUFX4_29/Y AOI21X1_191/B BUFX4_207/Y gnd AOI21X1_192/A vdd AOI21X1
XAOI21X1_180 AND2X2_24/Y BUFX4_57/Y AOI21X1_180/C gnd OAI21X1_517/A vdd AOI21X1
XNAND3X1_173 OR2X2_8/A OR2X2_8/B BUFX4_111/Y gnd XNOR2X1_8/A vdd NAND3X1
XNAND3X1_184 AOI21X1_43/A NAND2X1_145/Y NAND2X1_144/B gnd NAND3X1_185/C vdd NAND3X1
XFILL_31_5_1 gnd vdd FILL
XFILL_30_0_0 gnd vdd FILL
XNAND3X1_151 INVX8_10/Y OAI21X1_248/Y NAND3X1_151/C gnd NAND3X1_151/Y vdd NAND3X1
XNAND3X1_140 INVX1_82/Y NAND3X1_140/B NAND3X1_124/Y gnd NAND3X1_140/Y vdd NAND3X1
XNAND3X1_162 INVX4_4/Y NAND3X1_162/B NAND3X1_161/Y gnd NAND3X1_162/Y vdd NAND3X1
XNAND3X1_195 OR2X2_10/Y AOI21X1_34/B OAI21X1_277/C gnd AOI21X1_49/A vdd NAND3X1
XFILL_22_5_1 gnd vdd FILL
XOAI21X1_358 INVX2_52/Y BUFX4_162/Y OAI21X1_587/C gnd OAI21X1_358/Y vdd OAI21X1
XFILL_21_0_0 gnd vdd FILL
XOAI21X1_369 INVX2_120/Y BUFX4_161/Y NAND2X1_222/Y gnd AOI21X1_117/B vdd OAI21X1
XOAI21X1_303 AOI21X1_49/Y AOI21X1_50/Y INVX1_109/Y gnd INVX1_126/A vdd OAI21X1
XOAI21X1_336 BUFX4_223/Y BUFX4_234/Y DFFSR_239/Q gnd OAI21X1_336/Y vdd OAI21X1
XOAI21X1_325 OAI21X1_325/A OAI21X1_324/Y OAI21X1_325/C gnd DFFSR_242/D vdd OAI21X1
XOAI21X1_347 NOR2X1_209/Y MUX2X1_3/B BUFX4_55/Y gnd AOI21X1_109/C vdd OAI21X1
XOAI21X1_314 NAND2X1_197/Y NAND2X1_198/Y INVX2_164/A gnd OAI21X1_314/Y vdd OAI21X1
XDFFSR_182 INVX2_73/A CLKBUF1_13/Y DFFSR_137/R vdd DFFSR_182/D gnd vdd DFFSR
XNAND2X1_320 BUFX4_208/Y NAND2X1_320/B gnd OAI21X1_725/C vdd NAND2X1
XDFFSR_171 INVX2_129/A CLKBUF1_50/Y DFFSR_203/R vdd DFFSR_171/D gnd vdd DFFSR
XBUFX4_1 BUFX4_1/A gnd BUFX4_1/Y vdd BUFX4
XDFFSR_193 INVX1_58/A DFFSR_28/CLK DFFSR_130/R vdd DFFSR_193/D gnd vdd DFFSR
XDFFSR_160 INVX1_56/A CLKBUF1_33/Y DFFSR_167/R vdd DFFSR_160/D gnd vdd DFFSR
XNAND2X1_342 DFFSR_33/Q INVX4_5/Y gnd OAI21X1_791/C vdd NAND2X1
XFILL_29_1_0 gnd vdd FILL
XFILL_4_1_0 gnd vdd FILL
XNAND2X1_331 INVX2_126/A BUFX4_205/Y gnd NAND2X1_331/Y vdd NAND2X1
XFILL_5_6_1 gnd vdd FILL
XINVX4_1 wb_adr_i[2] gnd INVX4_1/Y vdd INVX4
XFILL_12_0_0 gnd vdd FILL
XFILL_13_5_1 gnd vdd FILL
XNAND3X1_4 BUFX4_14/Y NAND3X1_4/B BUFX4_22/Y gnd NAND3X1_4/Y vdd NAND3X1
XOAI21X1_133 BUFX4_93/Y BUFX4_103/Y DFFSR_7/Q gnd BUFX2_9/A vdd OAI21X1
XOAI21X1_188 OR2X2_8/B INVX2_46/Y INVX1_83/A gnd NOR2X1_55/B vdd OAI21X1
XOAI21X1_144 BUFX4_93/Y BUFX4_103/Y INVX1_10/A gnd BUFX2_20/A vdd OAI21X1
XOAI21X1_122 INVX2_37/Y BUFX4_85/Y OAI21X1_90/C gnd NAND3X1_65/B vdd OAI21X1
XOAI21X1_111 AND2X2_3/Y INVX2_31/Y NAND3X1_59/Y gnd DFFSR_47/D vdd OAI21X1
XAOI22X1_9 INVX2_88/A AOI22X1_7/B INVX8_5/Y INVX2_91/A gnd AOI22X1_9/Y vdd AOI22X1
XOAI21X1_100 INVX2_26/Y BUFX4_6/Y OAI21X1_69/C gnd NAND3X1_54/B vdd OAI21X1
XOAI21X1_166 NOR2X1_41/Y NOR2X1_42/Y NOR2X1_46/B gnd OAI21X1_167/C vdd OAI21X1
XOAI21X1_199 XOR2X1_2/Y INVX8_9/Y OAI21X1_199/C gnd BUFX4_194/A vdd OAI21X1
XOAI21X1_155 BUFX4_91/Y BUFX4_97/Y INVX1_5/A gnd BUFX2_31/A vdd OAI21X1
XOAI21X1_177 OR2X2_5/A OR2X2_5/B DFFSR_112/Q gnd AOI22X1_34/D vdd OAI21X1
XNAND2X1_150 NAND2X1_150/A NAND2X1_150/B gnd INVX1_113/A vdd NAND2X1
XNAND2X1_161 INVX2_159/Y BUFX4_178/Y gnd AOI22X1_42/A vdd NAND2X1
XNAND2X1_19 BUFX4_9/Y wb_dat_i[10] gnd OAI21X1_67/C vdd NAND2X1
XNAND2X1_172 INVX2_106/Y BUFX4_154/Y gnd AOI22X1_47/D vdd NAND2X1
XNAND2X1_194 INVX2_76/Y BUFX4_176/Y gnd AOI22X1_66/C vdd NAND2X1
XNAND2X1_183 INVX2_97/Y BUFX4_173/Y gnd AOI22X1_53/A vdd NAND2X1
XAOI22X1_17 BUFX4_21/Y INVX1_1/A DFFSR_204/Q INVX8_5/Y gnd NAND3X1_94/C vdd AOI22X1
XAOI22X1_28 INVX2_151/A BUFX4_127/Y BUFX4_21/Y INVX1_6/A gnd NAND3X1_99/A vdd AOI22X1
XAOI22X1_39 AOI22X1_39/A AOI22X1_39/B AOI22X1_39/C AOI22X1_39/D gnd AOI22X1_39/Y vdd
+ AOI22X1
XFILL_5_1 gnd vdd FILL
XBUFX2_60 DFFSR_89/Q gnd wb_dat_o[24] vdd BUFX2
XFILL_27_4_1 gnd vdd FILL
XFILL_2_4_1 gnd vdd FILL
XFILL_10_3_1 gnd vdd FILL
XAOI21X1_50 INVX8_13/Y INVX2_45/Y AOI21X1_50/C gnd AOI21X1_50/Y vdd AOI21X1
XAOI21X1_72 INVX2_100/Y BUFX4_172/Y INVX1_118/A gnd AOI21X1_72/Y vdd AOI21X1
XAOI21X1_94 INVX2_77/Y BUFX4_157/Y AOI21X1_71/C gnd AOI21X1_94/Y vdd AOI21X1
XAOI21X1_61 INVX2_162/Y BUFX4_157/Y AOI21X1_71/C gnd AOI21X1_61/Y vdd AOI21X1
XOAI21X1_1 INVX1_1/Y MUX2X1_8/S OAI21X1_1/C gnd OAI21X1_1/Y vdd OAI21X1
XAOI21X1_83 INVX2_165/Y BUFX4_158/Y AOI21X1_71/C gnd AOI21X1_83/Y vdd AOI21X1
XFILL_9_0_0 gnd vdd FILL
XFILL_18_4_1 gnd vdd FILL
XXOR2X1_4 OR2X2_10/A XOR2X1_4/B gnd XOR2X1_4/Y vdd XOR2X1
XMUX2X1_5 wb_dat_i[29] MUX2X1_5/B BUFX4_73/Y gnd MUX2X1_5/Y vdd MUX2X1
XCLKBUF1_6 CLKBUF1_6/A gnd CLKBUF1_6/Y vdd CLKBUF1
XBUFX4_111 DFFSR_42/Q gnd BUFX4_111/Y vdd BUFX4
XBUFX4_144 INVX8_7/Y gnd DFFSR_7/R vdd BUFX4
XBUFX4_100 BUFX4_98/A gnd INVX4_5/A vdd BUFX4
XBUFX4_122 INVX8_20/Y gnd BUFX4_122/Y vdd BUFX4
XNOR2X1_215 OR2X2_12/B INVX8_14/Y gnd NOR2X1_215/Y vdd NOR2X1
XNOR2X1_204 INVX8_14/Y INVX1_123/Y gnd NOR2X1_204/Y vdd NOR2X1
XBUFX4_133 INVX8_24/Y gnd DFFSR_130/R vdd BUFX4
XBUFX4_166 INVX8_19/Y gnd BUFX4_166/Y vdd BUFX4
XBUFX4_155 BUFX4_154/A gnd BUFX4_155/Y vdd BUFX4
XBUFX4_177 BUFX4_172/A gnd BUFX4_177/Y vdd BUFX4
XBUFX4_188 BUFX4_185/A gnd BUFX4_188/Y vdd BUFX4
XFILL_33_2_1 gnd vdd FILL
XFILL_24_3 gnd vdd FILL
XNOR2X1_248 INVX4_7/Y NOR2X1_262/B gnd NOR2X1_248/Y vdd NOR2X1
XNOR2X1_226 NOR2X1_245/B OR2X2_12/A gnd NOR2X1_226/Y vdd NOR2X1
XBUFX4_199 BUFX4_200/A gnd BUFX4_199/Y vdd BUFX4
XNOR2X1_237 INVX2_110/A BUFX4_35/Y gnd NOR2X1_237/Y vdd NOR2X1
XNOR2X1_259 INVX2_72/A BUFX4_38/Y gnd NOR2X1_259/Y vdd NOR2X1
XFILL_24_2_1 gnd vdd FILL
XINVX8_8 wb_rst_i gnd INVX8_8/Y vdd INVX8
XBUFX4_28 BUFX4_32/A gnd BUFX4_28/Y vdd BUFX4
XBUFX4_39 BUFX4_36/A gnd BUFX4_39/Y vdd BUFX4
XFILL_7_3_1 gnd vdd FILL
XBUFX4_17 BUFX4_19/A gnd AND2X2_1/B vdd BUFX4
XFILL_15_2_1 gnd vdd FILL
XINVX2_100 DFFSR_132/Q gnd INVX2_100/Y vdd INVX2
XINVX2_144 INVX1_29/A gnd INVX2_144/Y vdd INVX2
XINVX2_133 INVX1_45/A gnd INVX2_133/Y vdd INVX2
XINVX2_122 INVX1_62/A gnd INVX2_122/Y vdd INVX2
XINVX2_111 INVX1_54/A gnd INVX2_111/Y vdd INVX2
XINVX2_155 INVX1_58/A gnd INVX2_155/Y vdd INVX2
XOAI21X1_529 AND2X2_26/Y INVX2_157/Y BUFX4_169/Y gnd AOI21X1_183/C vdd OAI21X1
XOAI21X1_507 BUFX4_57/Y AOI21X1_176/B OAI21X1_507/C gnd AOI21X1_177/B vdd OAI21X1
XOAI21X1_518 BUFX4_203/Y BUFX4_30/Y INVX2_98/A gnd OAI21X1_522/C vdd OAI21X1
XAOI21X1_170 INVX2_101/Y AOI21X1_170/B BUFX4_230/Y gnd OAI21X1_491/C vdd AOI21X1
XAOI21X1_192 AOI21X1_192/A OAI21X1_562/Y NOR2X1_267/Y gnd DFFSR_177/D vdd AOI21X1
XAOI21X1_181 NOR2X1_260/Y BUFX4_57/Y AOI21X1_181/C gnd OAI21X1_522/A vdd AOI21X1
XNAND3X1_174 BUFX4_111/Y AND2X2_9/Y AND2X2_18/Y gnd NOR2X1_177/B vdd NAND3X1
XNAND3X1_185 NOR2X1_179/Y OR2X2_11/Y NAND3X1_185/C gnd NAND3X1_191/B vdd NAND3X1
XFILL_30_0_1 gnd vdd FILL
XNAND3X1_196 INVX1_106/Y AND2X2_21/Y NAND3X1_191/Y gnd AOI21X1_69/C vdd NAND3X1
XNAND3X1_163 BUFX4_239/Y NAND3X1_163/B OAI21X1_262/Y gnd NAND3X1_165/B vdd NAND3X1
XNAND3X1_130 BUFX4_237/Y NAND3X1_130/B NAND3X1_130/C gnd NAND3X1_131/C vdd NAND3X1
XNAND3X1_152 BUFX4_237/Y NAND3X1_152/B NAND3X1_152/C gnd NAND3X1_153/C vdd NAND3X1
XNAND3X1_141 INVX8_10/Y OAI21X1_236/Y OAI21X1_237/Y gnd NAND3X1_141/Y vdd NAND3X1
XDFFSR_150 INVX1_31/A CLKBUF1_4/A DFFSR_137/R vdd DFFSR_150/D gnd vdd DFFSR
XOAI21X1_359 BUFX4_52/Y OAI21X1_358/Y BUFX4_241/Y gnd OAI21X1_359/Y vdd OAI21X1
XFILL_21_0_1 gnd vdd FILL
XOAI21X1_304 DFFSR_199/Q BUFX4_174/Y AOI21X1_88/Y gnd OAI21X1_304/Y vdd OAI21X1
XOAI21X1_337 NOR2X1_207/Y INVX2_108/Y BUFX4_53/Y gnd OAI21X1_337/Y vdd OAI21X1
XOAI21X1_326 BUFX4_223/Y BUFX4_234/Y INVX2_150/A gnd OAI21X1_330/C vdd OAI21X1
XOAI21X1_348 MUX2X1_3/B MUX2X1_8/S OAI21X1_458/C gnd OAI21X1_348/Y vdd OAI21X1
XOAI21X1_315 NAND2X1_199/Y NAND2X1_200/Y NOR2X1_191/Y gnd OAI21X1_315/Y vdd OAI21X1
XDFFSR_161 INVX1_57/A DFFSR_56/CLK DFFSR_130/R vdd DFFSR_161/D gnd vdd DFFSR
XNAND2X1_343 INVX2_42/Y INVX4_11/Y gnd OAI21X1_795/C vdd NAND2X1
XDFFSR_183 INVX1_33/A CLKBUF1_11/Y DFFSR_198/R vdd DFFSR_183/D gnd vdd DFFSR
XNAND2X1_332 INVX4_7/A AND2X2_32/A gnd NAND2X1_332/Y vdd NAND2X1
XNAND2X1_321 INVX8_23/A INVX1_151/Y gnd NOR2X1_321/A vdd NAND2X1
XDFFSR_194 INVX2_63/A CLKBUF1_34/A DFFSR_194/R vdd DFFSR_194/D gnd vdd DFFSR
XDFFSR_172 DFFSR_172/Q CLKBUF1_45/Y DFFSR_167/R vdd DFFSR_172/D gnd vdd DFFSR
XBUFX4_2 BUFX4_1/A gnd BUFX4_2/Y vdd BUFX4
XNAND2X1_310 INVX1_157/A BUFX4_62/Y gnd AOI22X1_83/C vdd NAND2X1
XFILL_29_1_1 gnd vdd FILL
XFILL_4_1_1 gnd vdd FILL
XINVX4_2 INVX4_2/A gnd INVX4_2/Y vdd INVX4
XFILL_12_0_1 gnd vdd FILL
XNAND3X1_5 BUFX4_14/Y NAND3X1_5/B BUFX4_23/Y gnd NAND3X1_5/Y vdd NAND3X1
XOAI21X1_112 INVX2_32/Y BUFX4_80/Y NAND2X1_26/Y gnd NAND3X1_60/B vdd OAI21X1
XOAI21X1_101 AND2X2_3/Y INVX2_26/Y NAND3X1_54/Y gnd DFFSR_58/D vdd OAI21X1
XOAI21X1_145 BUFX4_92/Y INVX4_5/A INVX1_11/A gnd BUFX2_21/A vdd OAI21X1
XOAI21X1_189 INVX1_85/Y NOR2X1_55/Y INVX2_18/A gnd OAI21X1_190/C vdd OAI21X1
XOAI21X1_134 BUFX4_95/Y BUFX4_102/Y DFFSR_8/Q gnd BUFX2_10/A vdd OAI21X1
XOAI21X1_123 AND2X2_3/Y INVX2_37/Y NAND3X1_65/Y gnd DFFSR_53/D vdd OAI21X1
XOAI21X1_167 INVX1_71/Y NOR2X1_46/B OAI21X1_167/C gnd DFFSR_104/D vdd OAI21X1
XOAI21X1_156 BUFX4_94/Y BUFX4_97/Y INVX1_6/A gnd BUFX2_32/A vdd OAI21X1
XOAI21X1_178 OR2X2_6/A OR2X2_6/B DFFSR_114/Q gnd AOI21X1_27/A vdd OAI21X1
XNAND2X1_140 INVX2_51/Y NAND2X1_138/B gnd AOI21X1_38/B vdd NAND2X1
XNAND2X1_151 INVX8_9/Y NAND2X1_151/B gnd OAI21X1_284/C vdd NAND2X1
XNAND2X1_173 INVX2_103/Y BUFX4_172/Y gnd AOI22X1_48/A vdd NAND2X1
XNAND2X1_195 INVX2_54/Y BUFX4_176/Y gnd AOI22X1_67/B vdd NAND2X1
XNAND2X1_162 INVX2_163/Y BUFX4_178/Y gnd AOI22X1_43/A vdd NAND2X1
XNAND2X1_184 INVX2_98/Y BUFX4_153/Y gnd AOI22X1_53/D vdd NAND2X1
XAOI22X1_29 INVX2_64/A BUFX4_124/Y INVX8_5/Y INVX2_66/A gnd AOI22X1_29/Y vdd AOI22X1
XAOI22X1_18 DFFSR_172/Q BUFX4_127/Y INVX8_6/Y INVX2_165/A gnd NAND3X1_94/A vdd AOI22X1
XOAI21X1_690 INVX2_100/Y BUFX4_160/Y NAND2X1_229/Y gnd NAND2X1_304/B vdd OAI21X1
XFILL_5_2 gnd vdd FILL
XBUFX2_50 DFFSR_79/Q gnd wb_dat_o[14] vdd BUFX2
XBUFX2_61 BUFX2_61/A gnd wb_dat_o[25] vdd BUFX2
XAOI21X1_40 AOI21X1_40/A AOI21X1_40/B INVX2_50/A gnd NOR2X1_179/B vdd AOI21X1
XAOI21X1_51 AOI21X1_37/Y AOI21X1_51/B INVX1_116/Y gnd AOI21X1_51/Y vdd AOI21X1
XAOI21X1_95 INVX2_75/Y BUFX4_154/Y AOI21X1_69/C gnd AOI22X1_66/D vdd AOI21X1
XAOI21X1_62 INVX2_161/Y BUFX4_176/Y INVX1_118/A gnd AOI22X1_43/C vdd AOI21X1
XOAI21X1_2 BUFX4_180/Y INVX1_1/Y OAI21X1_2/C gnd DFFSR_25/D vdd OAI21X1
XAOI21X1_84 INVX1_120/Y BUFX4_177/Y INVX1_118/A gnd AOI21X1_84/Y vdd AOI21X1
XFILL_9_0_1 gnd vdd FILL
XAOI21X1_73 INVX2_87/Y BUFX4_175/Y INVX1_117/A gnd AOI21X1_73/Y vdd AOI21X1
XFILL_20_6_0 gnd vdd FILL
XMUX2X1_6 wb_dat_i[28] INVX1_95/A MUX2X1_6/S gnd MUX2X1_6/Y vdd MUX2X1
XFILL_11_6_0 gnd vdd FILL
XCLKBUF1_7 CLKBUF1_7/A gnd CLKBUF1_7/Y vdd CLKBUF1
XBUFX4_101 BUFX4_98/A gnd BUFX4_101/Y vdd BUFX4
XBUFX4_145 INVX8_7/Y gnd DFFSR_2/R vdd BUFX4
XBUFX4_112 DFFSR_42/Q gnd BUFX4_112/Y vdd BUFX4
XBUFX4_134 INVX8_24/Y gnd DFFSR_137/R vdd BUFX4
XBUFX4_178 BUFX4_172/A gnd BUFX4_178/Y vdd BUFX4
XNOR2X1_249 BUFX4_150/Y OR2X2_12/B gnd INVX1_136/A vdd NOR2X1
XNOR2X1_216 OR2X2_13/B INVX8_14/Y gnd NOR2X1_216/Y vdd NOR2X1
XNOR2X1_227 INVX1_37/A BUFX4_244/Y gnd NOR2X1_227/Y vdd NOR2X1
XBUFX4_156 BUFX4_154/A gnd BUFX4_156/Y vdd BUFX4
XBUFX4_189 BUFX4_193/A gnd AOI21X1_7/B vdd BUFX4
XBUFX4_123 INVX8_20/Y gnd BUFX4_123/Y vdd BUFX4
XNOR2X1_238 BUFX4_148/Y NOR2X1_238/B gnd AND2X2_23/A vdd NOR2X1
XBUFX4_167 INVX8_19/Y gnd BUFX4_167/Y vdd BUFX4
XNOR2X1_205 INVX1_126/A INVX2_164/Y gnd INVX1_124/A vdd NOR2X1
XINVX8_9 INVX8_9/A gnd INVX8_9/Y vdd INVX8
XBUFX4_18 BUFX4_19/A gnd BUFX4_18/Y vdd BUFX4
XBUFX4_29 BUFX4_32/A gnd BUFX4_29/Y vdd BUFX4
XINVX2_101 DFFSR_196/Q gnd INVX2_101/Y vdd INVX2
XINVX2_145 INVX1_28/A gnd INVX2_145/Y vdd INVX2
XINVX2_134 INVX2_134/A gnd INVX2_134/Y vdd INVX2
XINVX2_112 INVX1_52/A gnd INVX2_112/Y vdd INVX2
XINVX2_123 DFFSR_163/Q gnd INVX2_123/Y vdd INVX2
XINVX2_156 DFFSR_129/Q gnd INVX2_156/Y vdd INVX2
XFILL_34_5_0 gnd vdd FILL
XOAI21X1_508 INVX2_113/Y BUFX4_12/Y OAI21X1_621/C gnd OAI21X1_509/B vdd OAI21X1
XOAI21X1_519 NOR2X1_260/Y INVX2_98/Y BUFX4_167/Y gnd AOI21X1_181/C vdd OAI21X1
XFILL_25_5_0 gnd vdd FILL
XFILL_0_5_0 gnd vdd FILL
XAOI21X1_171 AOI21X1_171/A OAI21X1_491/Y NOR2X1_254/Y gnd DFFSR_196/D vdd AOI21X1
XAOI21X1_182 AND2X2_25/Y BUFX4_66/Y AOI21X1_182/C gnd AOI21X1_182/Y vdd AOI21X1
XAOI21X1_193 INVX2_82/Y NAND2X1_259/Y BUFX4_29/Y gnd OAI21X1_564/C vdd AOI21X1
XAOI21X1_160 NOR2X1_242/Y BUFX4_57/Y AOI21X1_160/C gnd OAI21X1_464/A vdd AOI21X1
XFILL_8_6_0 gnd vdd FILL
XFILL_16_5_0 gnd vdd FILL
XNAND3X1_175 AND2X2_9/Y AND2X2_18/Y AND2X2_19/Y gnd NAND2X1_138/B vdd NAND3X1
XNAND3X1_186 BUFX4_111/Y NOR2X1_176/A OR2X2_8/Y gnd AOI21X1_44/B vdd NAND3X1
XNAND3X1_197 AOI21X1_37/C OR2X2_11/Y NAND3X1_185/C gnd AOI21X1_53/A vdd NAND3X1
XNAND3X1_120 BUFX4_239/Y NAND3X1_120/B OAI21X1_217/Y gnd NAND3X1_122/B vdd NAND3X1
XNAND3X1_164 INVX8_10/Y OAI21X1_263/Y OAI21X1_264/Y gnd NAND3X1_164/Y vdd NAND3X1
XNAND3X1_153 INVX4_4/A NAND3X1_151/Y NAND3X1_153/C gnd NAND3X1_153/Y vdd NAND3X1
XNAND3X1_131 INVX4_4/A NAND3X1_129/Y NAND3X1_131/C gnd NAND3X1_131/Y vdd NAND3X1
XNAND3X1_142 MUX2X1_1/S OAI21X1_238/Y OAI21X1_239/Y gnd NAND3X1_142/Y vdd NAND3X1
XOAI21X1_305 INVX1_33/A BUFX4_174/Y AOI21X1_89/Y gnd NAND3X1_204/B vdd OAI21X1
XDFFSR_151 INVX1_32/A CLKBUF1_19/Y DFFSR_151/R vdd DFFSR_151/D gnd vdd DFFSR
XDFFSR_184 INVX1_36/A CLKBUF1_6/Y DFFSR_198/R vdd DFFSR_184/D gnd vdd DFFSR
XOAI21X1_338 INVX2_108/Y BUFX4_72/Y OAI21X1_567/C gnd OAI21X1_338/Y vdd OAI21X1
XOAI21X1_349 BUFX4_55/Y OAI21X1_348/Y BUFX4_240/Y gnd OAI21X1_349/Y vdd OAI21X1
XDFFSR_173 DFFSR_173/Q CLKBUF1_42/Y DFFSR_194/R vdd DFFSR_173/D gnd vdd DFFSR
XDFFSR_140 INVX1_120/A CLKBUF1_2/Y DFFSR_174/R vdd DFFSR_140/D gnd vdd DFFSR
XOAI21X1_316 NOR2X1_188/Y INVX2_125/Y BUFX4_56/Y gnd AOI21X1_103/C vdd OAI21X1
XOAI21X1_327 NOR2X1_204/Y INVX2_150/Y BUFX4_53/Y gnd AOI21X1_105/C vdd OAI21X1
XBUFX4_3 BUFX4_1/A gnd BUFX4_3/Y vdd BUFX4
XDFFSR_162 INVX2_61/A CLKBUF1_28/Y DFFSR_130/R vdd DFFSR_162/D gnd vdd DFFSR
XNAND2X1_344 INVX2_49/A INVX4_5/Y gnd NAND2X1_344/Y vdd NAND2X1
XNAND2X1_322 BUFX4_211/Y NAND2X1_322/B gnd NAND2X1_322/Y vdd NAND2X1
XNAND2X1_300 INVX2_80/Y NAND2X1_299/Y gnd OAI21X1_684/C vdd NAND2X1
XNAND2X1_333 BUFX4_82/Y wb_dat_i[7] gnd OAI21X1_787/C vdd NAND2X1
XDFFSR_195 INVX1_63/A CLKBUF1_34/A DFFSR_167/R vdd DFFSR_195/D gnd vdd DFFSR
XNAND2X1_311 INVX8_23/A INVX1_146/A gnd OAI21X1_704/B vdd NAND2X1
XINVX4_3 INVX4_3/A gnd INVX4_3/Y vdd INVX4
XFILL_31_3_0 gnd vdd FILL
XNAND3X1_6 BUFX4_14/Y NAND3X1_6/B BUFX4_22/Y gnd OAI21X1_8/C vdd NAND3X1
XOAI21X1_146 BUFX4_92/Y INVX4_5/A DFFSR_20/Q gnd BUFX2_22/A vdd OAI21X1
XOAI21X1_113 AND2X2_3/Y INVX2_32/Y NAND3X1_60/Y gnd DFFSR_48/D vdd OAI21X1
XOAI21X1_124 INVX2_38/Y BUFX4_86/Y OAI21X1_92/C gnd NAND3X1_66/B vdd OAI21X1
XFILL_22_3_0 gnd vdd FILL
XOAI21X1_135 BUFX4_95/Y BUFX4_102/Y INVX2_1/A gnd BUFX2_11/A vdd OAI21X1
XOAI21X1_102 INVX2_27/Y BUFX4_7/Y OAI21X1_71/C gnd NAND3X1_55/B vdd OAI21X1
XOAI21X1_157 BUFX4_94/Y BUFX4_97/Y INVX1_7/A gnd BUFX2_33/A vdd OAI21X1
XOAI21X1_168 BUFX4_4/Y XNOR2X1_1/Y NAND2X1_92/Y gnd DFFSR_105/D vdd OAI21X1
XOAI21X1_179 OR2X2_6/A INVX1_78/Y NOR2X1_46/B gnd OAI21X1_179/Y vdd OAI21X1
XNAND2X1_141 NAND2X1_141/A AOI21X1_39/A gnd AOI21X1_37/C vdd NAND2X1
XNAND2X1_130 INVX4_3/Y NOR2X1_180/B gnd AOI21X1_43/A vdd NAND2X1
XNAND2X1_152 INVX2_144/Y BUFX4_172/Y gnd AOI22X1_37/A vdd NAND2X1
XNAND2X1_174 INVX2_101/Y BUFX4_154/Y gnd AOI22X1_48/D vdd NAND2X1
XNAND2X1_196 INVX2_58/Y BUFX4_178/Y gnd AOI22X1_67/C vdd NAND2X1
XNAND2X1_163 INVX2_160/Y BUFX4_157/Y gnd AOI22X1_43/D vdd NAND2X1
XNAND2X1_185 INVX2_121/Y BUFX4_175/Y gnd AOI22X1_55/B vdd NAND2X1
XFILL_5_4_0 gnd vdd FILL
XFILL_13_3_0 gnd vdd FILL
XOAI21X1_691 INVX1_153/Y DFFSR_132/Q BUFX4_113/Y gnd OAI21X1_691/Y vdd OAI21X1
XOAI21X1_680 BUFX4_96/Y INVX8_18/Y NOR2X1_278/Y gnd INVX1_151/A vdd OAI21X1
XAOI22X1_19 DFFSR_173/Q BUFX4_124/Y INVX8_5/Y DFFSR_205/Q gnd NAND3X1_95/B vdd AOI22X1
XFILL_5_3 gnd vdd FILL
XBUFX2_40 BUFX2_40/A gnd wb_dat_o[4] vdd BUFX2
XBUFX2_62 BUFX2_62/A gnd wb_dat_o[26] vdd BUFX2
XBUFX2_51 BUFX2_51/A gnd wb_dat_o[15] vdd BUFX2
XAOI21X1_41 INVX1_105/Y AOI21X1_41/B INVX8_9/Y gnd AOI22X1_36/C vdd AOI21X1
XAOI21X1_52 INVX2_145/Y BUFX4_154/Y AOI21X1_69/C gnd AOI22X1_37/B vdd AOI21X1
XAOI21X1_30 AOI21X1_30/A AOI21X1_30/B BUFX4_41/Y gnd AOI21X1_30/Y vdd AOI21X1
XAOI21X1_96 INVX2_80/Y BUFX4_176/Y INVX1_118/A gnd AOI21X1_96/Y vdd AOI21X1
XOAI21X1_3 INVX1_2/Y BUFX4_71/Y OAI21X1_3/C gnd NAND3X1_4/B vdd OAI21X1
XAOI21X1_74 INVX1_95/Y BUFX4_177/Y INVX1_118/A gnd AOI21X1_74/Y vdd AOI21X1
XAOI21X1_63 MUX2X1_3/A BUFX4_153/Y AOI21X1_69/C gnd AOI21X1_63/Y vdd AOI21X1
XAOI21X1_85 AOI21X1_85/A AOI21X1_85/B INVX1_126/A gnd NOR3X1_3/C vdd AOI21X1
XFILL_20_6_1 gnd vdd FILL
XFILL_27_2_0 gnd vdd FILL
XFILL_2_2_0 gnd vdd FILL
XMUX2X1_7 wb_dat_i[27] INVX1_96/A MUX2X1_7/S gnd MUX2X1_7/Y vdd MUX2X1
XFILL_11_6_1 gnd vdd FILL
XCLKBUF1_8 CLKBUF1_8/A gnd CLKBUF1_8/Y vdd CLKBUF1
XFILL_10_1_0 gnd vdd FILL
XBUFX4_102 BUFX4_98/A gnd BUFX4_102/Y vdd BUFX4
XBUFX4_146 INVX8_7/Y gnd DFFSR_88/R vdd BUFX4
XBUFX4_179 AND2X2_1/Y gnd BUFX4_179/Y vdd BUFX4
XBUFX4_113 INVX8_21/Y gnd BUFX4_113/Y vdd BUFX4
XNOR2X1_217 AOI22X1_2/C BUFX4_241/Y gnd NOR2X1_217/Y vdd NOR2X1
XBUFX4_157 BUFX4_154/A gnd BUFX4_157/Y vdd BUFX4
XBUFX4_135 INVX8_24/Y gnd DFFSR_198/R vdd BUFX4
XFILL_18_2_0 gnd vdd FILL
XNOR2X1_228 INVX1_128/A OR2X2_12/A gnd NOR2X1_228/Y vdd NOR2X1
XBUFX4_124 NOR3X1_1/Y gnd BUFX4_124/Y vdd BUFX4
XBUFX4_168 INVX8_19/Y gnd BUFX4_168/Y vdd BUFX4
XNOR2X1_206 INVX8_14/Y INVX1_124/Y gnd NOR2X1_206/Y vdd NOR2X1
XNOR2X1_239 INVX8_15/A NOR2X1_239/B gnd AND2X2_24/A vdd NOR2X1
XBUFX4_19 BUFX4_19/A gnd BUFX4_19/Y vdd BUFX4
XINVX2_102 AOI22X1_2/C gnd INVX2_102/Y vdd INVX2
XINVX2_146 INVX2_146/A gnd INVX2_146/Y vdd INVX2
XINVX2_157 INVX1_39/A gnd INVX2_157/Y vdd INVX2
XINVX2_135 DFFSR_123/Q gnd INVX2_135/Y vdd INVX2
XINVX2_124 INVX1_63/A gnd INVX2_124/Y vdd INVX2
XINVX2_113 INVX1_53/A gnd INVX2_113/Y vdd INVX2
XFILL_34_5_1 gnd vdd FILL
XFILL_33_0_0 gnd vdd FILL
XOAI21X1_509 BUFX4_222/Y OAI21X1_509/B BUFX4_49/Y gnd AOI21X1_177/A vdd OAI21X1
XFILL_15_1 gnd vdd FILL
XFILL_25_5_1 gnd vdd FILL
XFILL_0_5_1 gnd vdd FILL
XFILL_24_0_0 gnd vdd FILL
XAOI21X1_150 INVX2_66/Y NAND2X1_248/Y BUFX4_234/Y gnd OAI21X1_435/C vdd AOI21X1
XAOI21X1_161 INVX2_55/Y OAI21X1_465/B BUFX4_230/Y gnd AOI21X1_161/Y vdd AOI21X1
XAOI21X1_183 AND2X2_26/Y BUFX4_60/Y AOI21X1_183/C gnd OAI21X1_532/A vdd AOI21X1
XAOI21X1_194 BUFX4_29/Y AOI21X1_194/B BUFX4_207/Y gnd AOI21X1_195/A vdd AOI21X1
XAOI21X1_172 INVX2_63/Y AOI21X1_172/B BUFX4_231/Y gnd OAI21X1_494/C vdd AOI21X1
XFILL_7_1_0 gnd vdd FILL
XFILL_8_6_1 gnd vdd FILL
XNAND3X1_121 INVX8_10/Y NAND3X1_121/B NAND3X1_121/C gnd NAND3X1_121/Y vdd NAND3X1
XNAND3X1_110 INVX8_10/Y NAND3X1_110/B NAND3X1_110/C gnd NAND3X1_110/Y vdd NAND3X1
XNAND3X1_132 INVX2_47/Y NAND3X1_128/Y NAND3X1_131/Y gnd NAND3X1_139/C vdd NAND3X1
XFILL_16_5_1 gnd vdd FILL
XFILL_15_0_0 gnd vdd FILL
XNAND3X1_176 INVX2_51/Y AND2X2_19/Y AOI21X1_36/B gnd AOI21X1_40/A vdd NAND3X1
XNAND3X1_198 BUFX4_245/Y INVX1_115/A NAND3X1_198/C gnd NAND3X1_198/Y vdd NAND3X1
XNAND3X1_187 INVX2_46/A AOI21X1_44/A AOI21X1_44/B gnd OAI21X1_277/C vdd NAND3X1
XNAND3X1_165 INVX4_4/A NAND3X1_165/B NAND3X1_164/Y gnd NAND3X1_166/C vdd NAND3X1
XNAND3X1_154 INVX2_47/Y NAND3X1_153/Y NAND3X1_150/Y gnd NAND3X1_155/C vdd NAND3X1
XNAND3X1_143 INVX4_4/Y NAND3X1_141/Y NAND3X1_142/Y gnd NAND3X1_143/Y vdd NAND3X1
XOAI21X1_317 BUFX4_98/Y INVX8_11/Y BUFX4_37/Y gnd BUFX4_47/A vdd OAI21X1
XOAI21X1_306 INVX2_130/A BUFX4_174/Y AOI21X1_92/Y gnd NAND3X1_205/A vdd OAI21X1
XOAI21X1_328 INVX2_150/Y MUX2X1_7/S OAI21X1_328/C gnd OAI21X1_328/Y vdd OAI21X1
XDFFSR_196 DFFSR_196/Q DFFSR_1/CLK BUFX4_130/Y vdd DFFSR_196/D gnd vdd DFFSR
XDFFSR_152 INVX1_35/A CLKBUF1_13/Y DFFSR_151/R vdd DFFSR_152/D gnd vdd DFFSR
XDFFSR_185 INVX1_39/A CLKBUF1_1/Y DFFSR_198/R vdd DFFSR_185/D gnd vdd DFFSR
XOAI21X1_339 BUFX4_53/Y OAI21X1_338/Y BUFX4_242/Y gnd OAI21X1_339/Y vdd OAI21X1
XBUFX4_4 BUFX4_1/A gnd BUFX4_4/Y vdd BUFX4
XDFFSR_141 DFFSR_141/Q CLKBUF1_52/Y DFFSR_174/R vdd DFFSR_141/D gnd vdd DFFSR
XDFFSR_174 INVX2_68/A CLKBUF1_39/Y DFFSR_174/R vdd DFFSR_174/D gnd vdd DFFSR
XDFFSR_130 INVX1_91/A CLKBUF1_34/Y DFFSR_130/R vdd DFFSR_130/D gnd vdd DFFSR
XDFFSR_163 DFFSR_163/Q DFFSR_28/CLK DFFSR_130/R vdd DFFSR_163/D gnd vdd DFFSR
XNAND2X1_345 NOR2X1_50/A INVX4_5/A gnd NAND2X1_345/Y vdd NAND2X1
XNAND2X1_323 INVX8_23/A NOR2X1_309/Y gnd INVX1_159/A vdd NAND2X1
XNAND2X1_301 BUFX4_206/Y OAI21X1_685/Y gnd NAND2X1_301/Y vdd NAND2X1
XNAND2X1_334 INVX1_162/A BUFX4_62/Y gnd AOI22X1_84/C vdd NAND2X1
XNAND2X1_312 BUFX4_210/Y NAND2X1_312/B gnd OAI21X1_706/C vdd NAND2X1
XINVX4_4 INVX4_4/A gnd INVX4_4/Y vdd INVX4
XFILL_31_3_1 gnd vdd FILL
XNAND3X1_7 BUFX4_14/Y NAND3X1_7/B BUFX4_22/Y gnd NAND3X1_7/Y vdd NAND3X1
XOAI21X1_147 BUFX4_92/Y INVX4_5/A INVX1_13/A gnd BUFX2_23/A vdd OAI21X1
XOAI21X1_114 INVX2_33/Y BUFX4_81/Y NAND2X1_27/Y gnd NAND3X1_61/B vdd OAI21X1
XOAI21X1_125 AND2X2_3/Y INVX2_38/Y NAND3X1_66/Y gnd DFFSR_54/D vdd OAI21X1
XFILL_22_3_1 gnd vdd FILL
XOAI21X1_136 BUFX4_91/Y BUFX4_102/Y INVX2_2/A gnd BUFX2_12/A vdd OAI21X1
XOAI21X1_103 AND2X2_3/Y INVX2_27/Y NAND3X1_55/Y gnd DFFSR_59/D vdd OAI21X1
XOAI21X1_169 NAND2X1_94/Y XNOR2X1_1/B DFFSR_106/Q gnd AND2X2_7/A vdd OAI21X1
XOAI21X1_158 BUFX4_91/Y BUFX4_97/Y INVX1_8/A gnd BUFX2_34/A vdd OAI21X1
XBUFX2_1 BUFX2_1/A gnd mosi_pad_o vdd BUFX2
XNAND2X1_142 INVX2_42/A NOR2X1_177/B gnd NAND2X1_143/B vdd NAND2X1
XNAND2X1_153 AOI21X1_43/Y AOI21X1_45/B gnd AOI21X1_51/B vdd NAND2X1
XNAND2X1_131 INVX1_104/Y INVX8_13/Y gnd AOI21X1_33/A vdd NAND2X1
XNAND2X1_175 AOI22X1_47/Y AOI22X1_48/Y gnd AOI22X1_50/B vdd NAND2X1
XNAND2X1_164 AOI22X1_42/Y AOI22X1_43/Y gnd AOI22X1_46/A vdd NAND2X1
XNAND2X1_186 INVX2_115/Y BUFX4_175/Y gnd AOI22X1_55/C vdd NAND2X1
XFILL_5_4_1 gnd vdd FILL
XNAND2X1_197 AOI22X1_69/Y AOI22X1_70/Y gnd NAND2X1_197/Y vdd NAND2X1
XNAND2X1_120 INVX2_99/Y INVX8_10/A gnd NAND2X1_120/Y vdd NAND2X1
XINVX2_1 INVX2_1/A gnd INVX2_1/Y vdd INVX2
XFILL_13_3_1 gnd vdd FILL
XOAI21X1_692 NOR2X1_313/Y OAI21X1_691/Y NAND2X1_304/Y gnd DFFSR_132/D vdd OAI21X1
XAOI21X1_1 DFFSR_116/Q AOI21X1_1/B AOI21X1_1/C gnd AOI21X1_1/Y vdd AOI21X1
XOAI21X1_670 OAI21X1_668/Y BUFX4_206/Y OAI21X1_670/C gnd DFFSR_138/D vdd OAI21X1
XOAI21X1_681 INVX1_151/A INVX8_22/Y INVX2_119/Y gnd OAI21X1_682/C vdd OAI21X1
XBUFX2_41 DFFSR_70/Q gnd wb_dat_o[5] vdd BUFX2
XBUFX2_52 DFFSR_81/Q gnd wb_dat_o[16] vdd BUFX2
XBUFX2_30 BUFX2_30/A gnd ss_pad_o[27] vdd BUFX2
XBUFX2_63 DFFSR_92/Q gnd wb_dat_o[27] vdd BUFX2
XAOI21X1_53 AOI21X1_53/A AOI21X1_53/B INVX8_9/Y gnd AOI21X1_53/Y vdd AOI21X1
XAOI21X1_42 INVX8_13/Y INVX1_90/A AOI21X1_42/C gnd INVX1_106/A vdd AOI21X1
XAOI21X1_86 INVX2_120/Y BUFX4_155/Y AOI21X1_71/C gnd AOI21X1_86/Y vdd AOI21X1
XAOI21X1_31 AOI21X1_31/A AOI21X1_31/B NOR2X1_76/B gnd AOI21X1_31/Y vdd AOI21X1
XAOI21X1_20 DFFSR_103/Q AND2X2_6/A AND2X2_5/Y gnd AOI21X1_20/Y vdd AOI21X1
XAOI21X1_64 MUX2X1_2/A BUFX4_173/Y INVX1_117/A gnd AOI21X1_64/Y vdd AOI21X1
XAOI21X1_75 INVX2_84/Y BUFX4_153/Y AOI21X1_69/C gnd AOI22X1_49/D vdd AOI21X1
XAOI21X1_97 INVX2_74/Y BUFX4_172/Y INVX1_117/A gnd AOI21X1_97/Y vdd AOI21X1
XOAI21X1_4 BUFX4_180/Y INVX1_2/Y NAND3X1_4/Y gnd DFFSR_26/D vdd OAI21X1
XFILL_27_2_1 gnd vdd FILL
XFILL_2_2_1 gnd vdd FILL
XMUX2X1_8 wb_dat_i[26] INVX1_93/A MUX2X1_8/S gnd MUX2X1_8/Y vdd MUX2X1
XFILL_10_1_1 gnd vdd FILL
XCLKBUF1_9 CLKBUF1_3/A gnd DFFSR_3/CLK vdd CLKBUF1
XBUFX4_103 BUFX4_98/A gnd BUFX4_103/Y vdd BUFX4
XBUFX4_114 INVX8_21/Y gnd BUFX4_114/Y vdd BUFX4
XBUFX4_125 NOR3X1_1/Y gnd AOI22X1_7/B vdd BUFX4
XBUFX4_136 INVX8_24/Y gnd DFFSR_174/R vdd BUFX4
XNOR2X1_229 INVX1_30/A BUFX4_241/Y gnd NOR2X1_229/Y vdd NOR2X1
XBUFX4_169 INVX8_19/Y gnd BUFX4_169/Y vdd BUFX4
XFILL_18_2_1 gnd vdd FILL
XBUFX4_147 INVX8_7/Y gnd DFFSR_95/R vdd BUFX4
XNOR2X1_207 INVX1_130/A INVX8_14/Y gnd NOR2X1_207/Y vdd NOR2X1
XNOR2X1_218 INVX1_61/A BUFX4_243/Y gnd NOR2X1_218/Y vdd NOR2X1
XBUFX4_158 BUFX4_154/A gnd BUFX4_158/Y vdd BUFX4
XINVX2_103 DFFSR_164/Q gnd INVX2_103/Y vdd INVX2
XINVX2_114 INVX1_34/A gnd INVX2_114/Y vdd INVX2
XINVX2_147 DFFSR_165/Q gnd INVX2_147/Y vdd INVX2
XINVX2_158 INVX1_40/A gnd INVX2_158/Y vdd INVX2
XINVX2_125 DFFSR_243/Q gnd INVX2_125/Y vdd INVX2
XINVX2_136 INVX1_49/A gnd MUX2X1_1/A vdd INVX2
XFILL_33_0_1 gnd vdd FILL
XFILL_15_2 gnd vdd FILL
XFILL_24_0_1 gnd vdd FILL
XAOI21X1_162 OAI21X1_467/Y OAI21X1_465/Y NOR2X1_244/Y gnd DFFSR_202/D vdd AOI21X1
XAOI21X1_184 NOR2X1_261/Y BUFX4_60/Y AOI21X1_184/C gnd OAI21X1_537/A vdd AOI21X1
XAOI21X1_140 NOR2X1_228/Y BUFX4_59/Y AOI21X1_140/C gnd OAI21X1_427/A vdd AOI21X1
XAOI21X1_151 AOI21X1_151/A AOI21X1_151/B NOR2X1_232/Y gnd DFFSR_210/D vdd AOI21X1
XAOI21X1_173 AOI21X1_173/A AOI21X1_173/B NOR2X1_255/Y gnd DFFSR_194/D vdd AOI21X1
XAOI21X1_195 AOI21X1_195/A AOI21X1_195/B NOR2X1_269/Y gnd DFFSR_176/D vdd AOI21X1
XFILL_7_1_1 gnd vdd FILL
XNAND3X1_111 BUFX4_239/Y OAI21X1_206/Y OAI21X1_207/Y gnd NAND3X1_112/C vdd NAND3X1
XNAND3X1_122 INVX4_4/A NAND3X1_122/B NAND3X1_121/Y gnd NAND3X1_123/C vdd NAND3X1
XNAND3X1_166 INVX2_47/Y NAND3X1_162/Y NAND3X1_166/C gnd NAND3X1_166/Y vdd NAND3X1
XNAND3X1_144 BUFX4_237/Y OAI21X1_240/Y NAND3X1_144/C gnd NAND3X1_146/B vdd NAND3X1
XFILL_15_0_1 gnd vdd FILL
XNAND3X1_100 NAND2X1_74/Y AOI22X1_29/Y AOI22X1_30/Y gnd DFFSR_95/D vdd NAND3X1
XNAND3X1_155 INVX1_84/Y NAND3X1_155/B NAND3X1_155/C gnd NAND3X1_155/Y vdd NAND3X1
XNAND3X1_133 INVX4_4/Y OAI21X1_229/Y OAI21X1_232/Y gnd NAND3X1_133/Y vdd NAND3X1
XNAND3X1_177 INVX2_50/A AOI21X1_40/A AOI21X1_40/B gnd NAND2X1_141/A vdd NAND3X1
XNAND3X1_188 INVX4_3/A OAI21X1_272/Y NOR2X1_177/B gnd NAND2X1_148/A vdd NAND3X1
XNAND3X1_199 INVX1_99/A OAI21X1_287/Y NAND3X1_198/Y gnd OAI21X1_293/C vdd NAND3X1
XOAI21X1_307 INVX2_134/A BUFX4_174/Y AOI21X1_93/Y gnd NAND3X1_205/B vdd OAI21X1
XOAI21X1_329 BUFX4_53/Y OAI21X1_328/Y BUFX4_242/Y gnd OAI21X1_329/Y vdd OAI21X1
XOAI21X1_318 INVX2_125/Y BUFX4_71/Y OAI21X1_738/C gnd OAI21X1_318/Y vdd OAI21X1
XDFFSR_164 DFFSR_164/Q CLKBUF1_6/A BUFX4_130/Y vdd DFFSR_164/D gnd vdd DFFSR
XDFFSR_153 INVX1_38/A CLKBUF1_12/Y DFFSR_137/R vdd DFFSR_153/D gnd vdd DFFSR
XNAND2X1_302 BUFX4_211/Y NAND2X1_302/B gnd OAI21X1_689/C vdd NAND2X1
XDFFSR_197 AOI22X1_3/D CLKBUF1_13/Y DFFSR_137/R vdd DFFSR_197/D gnd vdd DFFSR
XDFFSR_186 INVX1_42/A DFFSR_36/CLK DFFSR_198/R vdd DFFSR_186/D gnd vdd DFFSR
XDFFSR_120 INVX2_94/A CLKBUF1_12/A DFFSR_151/R vdd DFFSR_120/D gnd vdd DFFSR
XDFFSR_175 INVX2_109/A CLKBUF1_33/Y DFFSR_194/R vdd DFFSR_175/D gnd vdd DFFSR
XDFFSR_142 INVX1_93/A CLKBUF1_45/Y DFFSR_174/R vdd DFFSR_142/D gnd vdd DFFSR
XDFFSR_131 INVX1_98/A DFFSR_26/CLK DFFSR_130/R vdd DFFSR_131/D gnd vdd DFFSR
XBUFX4_5 wb_sel_i[1] gnd BUFX4_5/Y vdd BUFX4
XNAND2X1_346 INVX4_3/Y INVX4_2/Y gnd NOR2X1_347/A vdd NAND2X1
XNAND2X1_324 BUFX4_204/Y OAI21X1_729/Y gnd NAND2X1_324/Y vdd NAND2X1
XNAND2X1_335 INVX4_10/A AND2X2_31/A gnd AOI21X1_258/B vdd NAND2X1
XNAND2X1_313 BUFX4_210/Y NAND2X1_313/B gnd OAI21X1_710/C vdd NAND2X1
XINVX4_5 INVX4_5/A gnd INVX4_5/Y vdd INVX4
XNAND3X1_8 BUFX4_14/Y NAND3X1_8/B BUFX4_22/Y gnd NAND3X1_8/Y vdd NAND3X1
XOAI21X1_148 BUFX4_92/Y INVX4_5/A DFFSR_22/Q gnd BUFX2_24/A vdd OAI21X1
XOAI21X1_115 AND2X2_3/Y INVX2_33/Y NAND3X1_61/Y gnd DFFSR_49/D vdd OAI21X1
XOAI21X1_126 INVX4_1/Y NAND2X1_34/Y NOR2X1_19/B gnd BUFX4_193/A vdd OAI21X1
XOAI21X1_104 INVX2_28/Y BUFX4_8/Y OAI21X1_73/C gnd NAND3X1_56/B vdd OAI21X1
XOAI21X1_137 BUFX4_91/Y NOR2X1_1/A INVX2_3/A gnd BUFX2_13/A vdd OAI21X1
XOAI21X1_159 NAND2X1_85/B OR2X2_3/Y NAND2X1_85/Y gnd DFFSR_99/D vdd OAI21X1
XNAND2X1_143 NAND3X1_180/Y NAND2X1_143/B gnd OR2X2_11/A vdd NAND2X1
XNAND2X1_132 INVX4_2/A XNOR2X1_8/Y gnd NAND2X1_136/A vdd NAND2X1
XNAND2X1_121 INVX2_100/Y BUFX4_217/Y gnd NAND3X1_134/C vdd NAND2X1
XNAND2X1_110 INVX1_87/A XOR2X1_2/B gnd NAND2X1_110/Y vdd NAND2X1
XBUFX2_2 BUFX2_2/A gnd sclk_pad_o vdd BUFX2
XNAND2X1_154 INVX2_147/Y BUFX4_172/Y gnd AOI22X1_38/B vdd NAND2X1
XNAND2X1_187 INVX2_129/Y BUFX4_174/Y gnd AOI22X1_56/B vdd NAND2X1
XNAND2X1_198 AOI22X1_71/Y AOI22X1_72/Y gnd NAND2X1_198/Y vdd NAND2X1
XNAND2X1_165 MUX2X1_1/A BUFX4_173/Y gnd AOI22X1_44/A vdd NAND2X1
XNAND2X1_176 INVX2_85/Y BUFX4_173/Y gnd AOI22X1_49/C vdd NAND2X1
XINVX2_2 INVX2_2/A gnd INVX2_2/Y vdd INVX2
XOAI21X1_671 BUFX4_58/Y NAND2X1_292/Y NAND2X1_293/Y gnd OAI21X1_673/A vdd OAI21X1
XAOI21X1_2 INVX1_99/A AOI21X1_2/B AOI21X1_2/C gnd AOI21X1_2/Y vdd AOI21X1
XOAI21X1_682 BUFX4_64/Y OAI21X1_682/B OAI21X1_682/C gnd OAI21X1_683/A vdd OAI21X1
XOAI21X1_660 MUX2X1_2/B BUFX4_70/Y OAI21X1_458/C gnd OAI21X1_660/Y vdd OAI21X1
XOAI21X1_693 INVX1_91/Y BUFX4_7/Y NAND2X1_231/Y gnd NAND2X1_306/B vdd OAI21X1
XXNOR2X1_10 XNOR2X1_8/Y INVX4_2/Y gnd XNOR2X1_10/Y vdd XNOR2X1
XBUFX2_53 BUFX2_53/A gnd wb_dat_o[17] vdd BUFX2
XBUFX2_42 BUFX2_42/A gnd wb_dat_o[6] vdd BUFX2
XFILL_32_6_0 gnd vdd FILL
XBUFX2_20 BUFX2_20/A gnd ss_pad_o[17] vdd BUFX2
XBUFX2_31 BUFX2_31/A gnd ss_pad_o[28] vdd BUFX2
XBUFX2_64 BUFX2_64/A gnd wb_dat_o[28] vdd BUFX2
XFILL_23_6_0 gnd vdd FILL
XAOI21X1_43 AOI21X1_43/A AOI21X1_43/B NOR2X1_180/Y gnd AOI21X1_43/Y vdd AOI21X1
XAOI21X1_54 AOI21X1_43/Y AOI21X1_45/B AOI21X1_54/C gnd AOI21X1_54/Y vdd AOI21X1
XAOI21X1_32 INVX1_17/A INVX2_53/Y BUFX4_245/Y gnd AOI21X1_32/Y vdd AOI21X1
XAOI21X1_98 INVX2_52/Y BUFX4_157/Y AOI21X1_71/C gnd AOI21X1_98/Y vdd AOI21X1
XAOI21X1_87 INVX2_114/Y BUFX4_156/Y AOI21X1_69/C gnd AOI22X1_55/D vdd AOI21X1
XAOI21X1_10 INVX2_138/A AOI21X1_7/B AOI21X1_10/C gnd NAND2X1_51/A vdd AOI21X1
XOAI21X1_5 INVX1_3/Y BUFX4_73/Y OAI21X1_5/C gnd NAND3X1_5/B vdd OAI21X1
XAOI21X1_21 NOR2X1_40/Y NOR2X1_27/Y OR2X2_1/A gnd NOR2X1_46/B vdd AOI21X1
XAOI21X1_65 MUX2X1_3/B BUFX4_153/Y AOI21X1_71/C gnd AOI21X1_65/Y vdd AOI21X1
XAOI21X1_76 INVX2_81/Y BUFX4_153/Y AOI21X1_71/C gnd AOI21X1_76/Y vdd AOI21X1
XFILL_14_6_0 gnd vdd FILL
XOAI22X1_40 OAI22X1_41/A OR2X2_1/Y NAND2X1_82/Y OAI22X1_40/D gnd DFFSR_97/D vdd OAI22X1
XOAI21X1_490 AOI21X1_169/Y OAI21X1_490/B OAI21X1_490/C gnd DFFSR_197/D vdd OAI21X1
XMUX2X1_9 wb_dat_i[11] INVX1_97/A BUFX4_10/Y gnd MUX2X1_9/Y vdd MUX2X1
XBUFX4_159 wb_sel_i[2] gnd NAND2X1_9/B vdd BUFX4
XBUFX4_126 NOR3X1_1/Y gnd AOI22X1_1/B vdd BUFX4
XBUFX4_115 INVX8_21/Y gnd BUFX4_115/Y vdd BUFX4
XBUFX4_137 INVX8_24/Y gnd DFFSR_194/R vdd BUFX4
XBUFX4_104 BUFX4_98/A gnd NOR2X1_1/A vdd BUFX4
XBUFX4_148 BUFX4_152/A gnd BUFX4_148/Y vdd BUFX4
XNOR2X1_208 NOR2X1_238/B INVX8_14/Y gnd NOR2X1_208/Y vdd NOR2X1
XNOR2X1_219 OR2X2_12/A INVX1_123/Y gnd NOR2X1_219/Y vdd NOR2X1
XFILL_20_4_0 gnd vdd FILL
XFILL_28_5_0 gnd vdd FILL
XFILL_3_5_0 gnd vdd FILL
XINVX2_104 INVX1_26/A gnd INVX2_104/Y vdd INVX2
XINVX2_115 INVX1_32/A gnd INVX2_115/Y vdd INVX2
XINVX2_137 DFFSR_173/Q gnd MUX2X1_1/B vdd INVX2
XINVX2_126 INVX2_126/A gnd INVX2_126/Y vdd INVX2
XFILL_11_4_0 gnd vdd FILL
XINVX2_159 INVX1_38/A gnd INVX2_159/Y vdd INVX2
XINVX2_148 AOI22X1_4/C gnd INVX2_148/Y vdd INVX2
XFILL_19_5_0 gnd vdd FILL
XAOI21X1_141 INVX2_75/Y OR2X2_12/Y BUFX4_151/Y gnd AOI21X1_141/Y vdd AOI21X1
XAOI21X1_185 NOR2X1_262/Y BUFX4_66/Y AOI21X1_185/C gnd AOI21X1_185/Y vdd AOI21X1
XAOI21X1_163 INVX2_160/Y AOI21X1_163/B BUFX4_230/Y gnd OAI21X1_468/C vdd AOI21X1
XAOI21X1_152 INVX2_152/Y OR2X2_14/Y BUFX4_234/Y gnd OAI21X1_439/C vdd AOI21X1
XAOI21X1_196 AND2X2_29/Y BUFX4_63/Y AOI21X1_196/C gnd OAI21X1_569/A vdd AOI21X1
XAOI21X1_130 BUFX4_148/Y OAI21X1_395/Y BUFX4_49/Y gnd AOI21X1_131/A vdd AOI21X1
XAOI21X1_174 NOR2X1_256/Y BUFX4_57/Y AOI21X1_174/C gnd AOI21X1_174/Y vdd AOI21X1
XNAND3X1_178 OR2X2_7/B AND2X2_19/Y AOI21X1_36/B gnd XNOR2X1_9/A vdd NAND3X1
XNAND3X1_189 INVX4_3/Y NAND2X1_129/A NAND2X1_129/B gnd NAND2X1_148/B vdd NAND3X1
XNAND3X1_134 BUFX4_184/Y NAND3X1_134/B NAND3X1_134/C gnd NAND3X1_135/B vdd NAND3X1
XNAND3X1_156 BUFX4_239/Y OAI21X1_253/Y NAND3X1_156/C gnd NAND3X1_158/B vdd NAND3X1
XNAND3X1_112 INVX4_4/A NAND3X1_110/Y NAND3X1_112/C gnd NAND3X1_116/B vdd NAND3X1
XNAND3X1_167 INVX1_84/A NAND3X1_159/Y NAND3X1_166/Y gnd NAND3X1_167/Y vdd NAND3X1
XNAND3X1_123 INVX2_47/A NAND3X1_119/Y NAND3X1_123/C gnd NAND3X1_124/C vdd NAND3X1
XNAND3X1_145 INVX8_10/Y OAI21X1_242/Y OAI21X1_243/Y gnd NAND3X1_145/Y vdd NAND3X1
XNAND3X1_101 NAND2X1_75/Y AOI22X1_31/Y AOI22X1_32/Y gnd DFFSR_96/D vdd NAND3X1
XFILL_34_3_0 gnd vdd FILL
XFILL_20_1 gnd vdd FILL
XDFFSR_132 DFFSR_132/Q CLKBUF1_27/Y DFFSR_165/R vdd DFFSR_132/D gnd vdd DFFSR
XDFFSR_121 DFFSR_121/Q DFFSR_1/CLK BUFX4_130/Y vdd DFFSR_121/D gnd vdd DFFSR
XOAI21X1_319 BUFX4_55/Y OAI21X1_318/Y BUFX4_240/Y gnd OAI21X1_319/Y vdd OAI21X1
XDFFSR_110 INVX1_75/A CLKBUF1_2/Y vdd BUFX4_89/Y DFFSR_110/D gnd vdd DFFSR
XDFFSR_143 INVX1_96/A DFFSR_98/CLK DFFSR_174/R vdd DFFSR_143/D gnd vdd DFFSR
XOAI21X1_308 NAND2X1_189/Y NAND2X1_190/Y INVX2_164/A gnd OAI21X1_308/Y vdd OAI21X1
XNAND2X1_325 INVX8_23/A NOR2X1_310/Y gnd INVX1_160/A vdd NAND2X1
XDFFSR_165 DFFSR_165/Q CLKBUF1_54/Y DFFSR_165/R vdd DFFSR_165/D gnd vdd DFFSR
XNAND2X1_303 INVX8_22/A NOR2X1_310/Y gnd INVX1_152/A vdd NAND2X1
XDFFSR_198 INVX2_79/A CLKBUF1_11/Y DFFSR_198/R vdd DFFSR_198/D gnd vdd DFFSR
XDFFSR_154 INVX1_41/A CLKBUF1_5/Y DFFSR_151/R vdd DFFSR_154/D gnd vdd DFFSR
XDFFSR_187 INVX2_134/A CLKBUF1_48/Y DFFSR_198/R vdd DFFSR_187/D gnd vdd DFFSR
XNAND2X1_314 INVX8_23/A INVX1_149/A gnd OAI21X1_712/B vdd NAND2X1
XNAND2X1_336 INVX1_45/A INVX8_21/A gnd NAND2X1_336/Y vdd NAND2X1
XDFFSR_176 INVX2_82/A CLKBUF1_32/Y DFFSR_194/R vdd DFFSR_176/D gnd vdd DFFSR
XBUFX4_6 wb_sel_i[1] gnd BUFX4_6/Y vdd BUFX4
XNAND2X1_347 INVX2_50/Y INVX2_49/Y gnd NOR2X1_347/B vdd NAND2X1
XFILL_25_3_0 gnd vdd FILL
XINVX4_6 INVX4_6/A gnd INVX4_6/Y vdd INVX4
XFILL_0_3_0 gnd vdd FILL
XFILL_8_4_0 gnd vdd FILL
XFILL_16_3_0 gnd vdd FILL
XNAND3X1_9 BUFX4_14/Y NAND3X1_9/B BUFX4_22/Y gnd NAND3X1_9/Y vdd NAND3X1
XBUFX2_3 BUFX2_3/A gnd ss_pad_o[0] vdd BUFX2
XOAI21X1_127 BUFX4_92/Y BUFX4_103/Y DFFSR_1/Q gnd BUFX2_3/A vdd OAI21X1
XOAI21X1_149 BUFX4_93/Y BUFX4_102/Y INVX1_15/A gnd BUFX2_25/A vdd OAI21X1
XOAI21X1_116 INVX2_34/Y BUFX4_82/Y NAND2X1_28/Y gnd NAND3X1_62/B vdd OAI21X1
XOAI21X1_138 BUFX4_95/Y BUFX4_102/Y INVX2_4/A gnd BUFX2_14/A vdd OAI21X1
XOAI21X1_105 AND2X2_3/Y INVX2_28/Y NAND3X1_56/Y gnd DFFSR_60/D vdd OAI21X1
XNAND2X1_133 OR2X2_8/A OR2X2_8/B gnd NOR2X1_176/A vdd NAND2X1
XNAND2X1_144 AOI21X1_43/A NAND2X1_144/B gnd OAI21X1_275/A vdd NAND2X1
XNAND2X1_122 INVX2_101/Y BUFX4_45/Y gnd NAND3X1_134/B vdd NAND2X1
XNAND2X1_155 AOI22X1_37/Y AOI22X1_38/Y gnd AOI22X1_41/A vdd NAND2X1
XNAND2X1_111 INVX2_52/Y BUFX4_42/Y gnd NAND2X1_111/Y vdd NAND2X1
XNAND2X1_177 INVX2_82/Y BUFX4_177/Y gnd AOI22X1_49/B vdd NAND2X1
XNAND2X1_100 INVX2_30/A BUFX4_3/Y gnd OAI21X1_180/C vdd NAND2X1
XNAND2X1_166 MUX2X1_4/A BUFX4_155/Y gnd AOI22X1_44/D vdd NAND2X1
XNAND2X1_188 INVX2_133/Y BUFX4_174/Y gnd AOI22X1_56/C vdd NAND2X1
XNAND2X1_199 AOI22X1_73/Y AOI22X1_74/Y gnd NAND2X1_199/Y vdd NAND2X1
XOAI21X1_650 BUFX4_121/Y OAI21X1_649/Y BUFX4_114/Y gnd OAI21X1_650/Y vdd OAI21X1
XINVX2_3 INVX2_3/A gnd INVX2_3/Y vdd INVX2
XOAI21X1_672 INVX2_161/Y BUFX4_162/Y NAND2X1_216/Y gnd OAI21X1_672/Y vdd OAI21X1
XAOI21X1_3 INVX2_74/A AOI21X1_2/B AOI21X1_3/C gnd AOI21X1_3/Y vdd AOI21X1
XOAI21X1_683 OAI21X1_683/A BUFX4_208/Y OAI21X1_683/C gnd DFFSR_135/D vdd OAI21X1
XOAI21X1_661 INVX1_147/A DFFSR_141/Q BUFX4_117/Y gnd OAI21X1_662/B vdd OAI21X1
XOAI21X1_694 INVX1_154/A INVX1_91/A BUFX4_117/Y gnd OAI21X1_695/B vdd OAI21X1
XXNOR2X1_11 XNOR2X1_10/Y AOI21X1_34/Y gnd XNOR2X1_11/Y vdd XNOR2X1
XINVX1_90 INVX1_90/A gnd INVX1_90/Y vdd INVX1
XBUFX2_10 BUFX2_10/A gnd ss_pad_o[7] vdd BUFX2
XBUFX2_54 DFFSR_83/Q gnd wb_dat_o[18] vdd BUFX2
XBUFX2_21 BUFX2_21/A gnd ss_pad_o[18] vdd BUFX2
XFILL_32_6_1 gnd vdd FILL
XFILL_31_1_0 gnd vdd FILL
XBUFX2_43 BUFX2_43/A gnd wb_dat_o[7] vdd BUFX2
XBUFX2_32 BUFX2_32/A gnd ss_pad_o[29] vdd BUFX2
XBUFX2_65 DFFSR_94/Q gnd wb_dat_o[29] vdd BUFX2
XNOR2X1_1 NOR2X1_1/A NOR2X1_1/B gnd BUFX4_19/A vdd NOR2X1
XFILL_23_6_1 gnd vdd FILL
XFILL_22_1_0 gnd vdd FILL
XAOI21X1_44 AOI21X1_44/A AOI21X1_44/B INVX2_46/A gnd AOI21X1_44/Y vdd AOI21X1
XAOI21X1_33 AOI21X1_33/A AOI21X1_33/B INVX2_46/Y gnd AOI21X1_33/Y vdd AOI21X1
XAOI21X1_55 INVX2_148/Y BUFX4_154/Y AOI21X1_71/C gnd AOI21X1_55/Y vdd AOI21X1
XAOI21X1_99 INVX2_57/Y BUFX4_157/Y AOI21X1_69/C gnd AOI21X1_99/Y vdd AOI21X1
XAOI21X1_77 INVX2_93/Y BUFX4_156/Y AOI21X1_69/C gnd AOI21X1_77/Y vdd AOI21X1
XAOI21X1_88 INVX2_119/Y BUFX4_175/Y INVX1_118/A gnd AOI21X1_88/Y vdd AOI21X1
XOAI21X1_6 BUFX4_180/Y INVX1_3/Y NAND3X1_5/Y gnd DFFSR_27/D vdd OAI21X1
XAOI21X1_22 DFFSR_107/Q AND2X2_7/B NOR2X1_40/Y gnd AOI21X1_22/Y vdd AOI21X1
XAOI21X1_66 MUX2X1_2/B BUFX4_173/Y INVX1_118/A gnd AOI21X1_66/Y vdd AOI21X1
XAOI21X1_11 INVX1_94/A BUFX4_190/Y AOI21X1_11/C gnd NAND2X1_53/A vdd AOI21X1
XFILL_5_2_0 gnd vdd FILL
XOAI22X1_30 BUFX4_76/Y INVX2_5/Y INVX1_55/Y INVX8_6/A gnd NOR2X1_16/A vdd OAI22X1
XFILL_13_1_0 gnd vdd FILL
XOAI22X1_41 OAI22X1_41/A NAND2X1_83/Y NAND2X1_82/Y OR2X2_1/Y gnd DFFSR_98/D vdd OAI22X1
XFILL_14_6_1 gnd vdd FILL
XOAI21X1_491 BUFX4_61/Y AOI21X1_170/B OAI21X1_491/C gnd OAI21X1_491/Y vdd OAI21X1
XOAI21X1_480 OAI21X1_480/A OAI21X1_480/B OAI21X1_475/Y gnd DFFSR_199/D vdd OAI21X1
XBUFX4_105 INVX8_4/Y gnd AND2X2_3/A vdd BUFX4
XBUFX4_138 INVX8_24/Y gnd DFFSR_236/R vdd BUFX4
XBUFX4_127 NOR3X1_1/Y gnd BUFX4_127/Y vdd BUFX4
XBUFX4_116 INVX8_21/Y gnd BUFX4_116/Y vdd BUFX4
XNOR2X1_209 NOR2X1_239/B INVX8_14/Y gnd NOR2X1_209/Y vdd NOR2X1
XBUFX4_149 BUFX4_152/A gnd INVX8_15/A vdd BUFX4
XFILL_20_4_1 gnd vdd FILL
XFILL_28_5_1 gnd vdd FILL
XFILL_27_0_0 gnd vdd FILL
XFILL_3_5_1 gnd vdd FILL
XFILL_2_0_0 gnd vdd FILL
XFILL_11_4_1 gnd vdd FILL
XINVX2_105 INVX1_27/A gnd INVX2_105/Y vdd INVX2
XINVX2_149 AOI22X1_3/D gnd INVX2_149/Y vdd INVX2
XINVX2_116 INVX1_33/A gnd INVX2_116/Y vdd INVX2
XINVX2_127 INVX2_127/A gnd INVX2_127/Y vdd INVX2
XINVX2_138 INVX2_138/A gnd MUX2X1_2/A vdd INVX2
XFILL_19_5_1 gnd vdd FILL
XFILL_18_0_0 gnd vdd FILL
XINVX1_160 INVX1_160/A gnd INVX1_160/Y vdd INVX1
XAOI21X1_142 BUFX4_151/Y OAI21X1_429/Y BUFX4_47/Y gnd AOI21X1_142/Y vdd AOI21X1
XAOI21X1_186 NOR2X1_263/Y BUFX4_61/Y AOI21X1_186/C gnd OAI21X1_547/A vdd AOI21X1
XAOI21X1_120 NOR2X1_216/Y BUFX4_66/Y OAI21X1_376/Y gnd AOI21X1_120/Y vdd AOI21X1
XAOI21X1_164 AOI21X1_164/A AOI21X1_164/B NOR2X1_246/Y gnd DFFSR_201/D vdd AOI21X1
XAOI21X1_153 OAI21X1_441/Y AOI21X1_153/B NOR2X1_233/Y gnd DFFSR_209/D vdd AOI21X1
XAOI21X1_197 NOR2X1_271/Y BUFX4_63/Y AOI21X1_197/C gnd OAI21X1_574/A vdd AOI21X1
XAOI21X1_131 AOI21X1_131/A AOI21X1_131/B NOR2X1_221/Y gnd DFFSR_223/D vdd AOI21X1
XAOI21X1_175 NOR2X1_257/Y BUFX4_57/Y OAI21X1_503/Y gnd OAI21X1_506/A vdd AOI21X1
XNAND3X1_179 INVX2_50/Y XNOR2X1_9/A AOI21X1_38/B gnd AOI21X1_39/A vdd NAND3X1
XNAND3X1_135 INVX8_10/Y NAND3X1_135/B OAI21X1_233/Y gnd NAND3X1_135/Y vdd NAND3X1
XNAND3X1_157 INVX8_10/Y NAND3X1_157/B NAND3X1_157/C gnd NAND3X1_157/Y vdd NAND3X1
XNAND3X1_168 INVX1_82/A NAND3X1_167/Y NAND3X1_155/Y gnd NAND3X1_169/C vdd NAND3X1
XNAND3X1_146 INVX4_4/A NAND3X1_146/B NAND3X1_145/Y gnd NAND3X1_146/Y vdd NAND3X1
XNAND3X1_124 INVX1_84/Y NAND3X1_124/B NAND3X1_124/C gnd NAND3X1_124/Y vdd NAND3X1
XNAND3X1_102 XOR2X1_1/A INVX1_65/Y AND2X2_5/A gnd NOR2X1_31/B vdd NAND3X1
XNAND3X1_113 BUFX4_238/Y OAI21X1_208/Y OAI21X1_209/Y gnd NAND3X1_113/Y vdd NAND3X1
XFILL_34_3_1 gnd vdd FILL
XFILL_20_2 gnd vdd FILL
XDFFSR_133 DFFSR_133/Q DFFSR_88/CLK DFFSR_137/R vdd DFFSR_133/D gnd vdd DFFSR
XDFFSR_166 INVX2_78/A DFFSR_1/CLK BUFX4_130/Y vdd DFFSR_166/D gnd vdd DFFSR
XDFFSR_122 INVX2_60/A CLKBUF1_13/Y DFFSR_151/R vdd DFFSR_122/D gnd vdd DFFSR
XDFFSR_155 INVX1_45/A DFFSR_5/CLK DFFSR_151/R vdd DFFSR_155/D gnd vdd DFFSR
XBUFX4_7 wb_sel_i[1] gnd BUFX4_7/Y vdd BUFX4
XDFFSR_144 INVX1_95/A DFFSR_99/CLK DFFSR_174/R vdd DFFSR_144/D gnd vdd DFFSR
XDFFSR_111 OR2X2_5/B CLKBUF1_52/Y vdd BUFX4_90/Y DFFSR_111/D gnd vdd DFFSR
XOAI21X1_309 NAND2X1_191/Y NAND2X1_192/Y NOR2X1_191/Y gnd OAI21X1_309/Y vdd OAI21X1
XDFFSR_100 XOR2X1_1/A CLKBUF1_35/Y vdd BUFX4_89/Y DFFSR_100/D gnd vdd DFFSR
XFILL_13_1 gnd vdd FILL
XNAND2X1_326 BUFX4_204/Y OAI21X1_732/Y gnd NAND2X1_326/Y vdd NAND2X1
XNAND2X1_304 BUFX4_204/Y NAND2X1_304/B gnd NAND2X1_304/Y vdd NAND2X1
XNAND2X1_315 BUFX4_208/Y NAND2X1_315/B gnd OAI21X1_714/C vdd NAND2X1
XDFFSR_199 DFFSR_199/Q CLKBUF1_6/Y DFFSR_198/R vdd DFFSR_199/D gnd vdd DFFSR
XDFFSR_177 INVX2_151/A CLKBUF1_26/Y DFFSR_174/R vdd DFFSR_177/D gnd vdd DFFSR
XNAND2X1_337 BUFX4_205/Y NAND2X1_337/B gnd OAI21X1_782/C vdd NAND2X1
XDFFSR_188 INVX2_98/A CLKBUF1_42/Y DFFSR_167/R vdd DFFSR_188/D gnd vdd DFFSR
XFILL_25_3_1 gnd vdd FILL
XFILL_0_3_1 gnd vdd FILL
XINVX4_7 INVX4_7/A gnd INVX4_7/Y vdd INVX4
XFILL_8_4_1 gnd vdd FILL
XFILL_16_3_1 gnd vdd FILL
XOAI21X1_128 BUFX4_92/Y BUFX4_103/Y DFFSR_2/Q gnd BUFX2_4/A vdd OAI21X1
XOAI21X1_117 AND2X2_3/Y INVX2_34/Y NAND3X1_62/Y gnd DFFSR_50/D vdd OAI21X1
XOAI21X1_106 INVX2_29/Y BUFX4_9/Y OAI21X1_45/C gnd NAND3X1_57/B vdd OAI21X1
XBUFX2_4 BUFX2_4/A gnd ss_pad_o[1] vdd BUFX2
XOAI21X1_139 BUFX4_95/Y BUFX4_102/Y INVX2_5/A gnd BUFX2_15/A vdd OAI21X1
XNAND2X1_145 AND2X2_20/B AND2X2_20/A gnd NAND2X1_145/Y vdd NAND2X1
XNAND2X1_134 BUFX4_111/Y INVX2_43/Y gnd NAND2X1_134/Y vdd NAND2X1
XNAND2X1_101 INVX2_43/Y NOR2X1_47/Y gnd NOR2X1_48/B vdd NAND2X1
XNAND2X1_112 OR2X2_9/B OR2X2_9/A gnd NAND3X1_108/B vdd NAND2X1
XNAND2X1_178 INVX2_92/Y BUFX4_178/Y gnd AOI22X1_51/A vdd NAND2X1
XNAND2X1_189 AOI22X1_58/Y AOI22X1_59/Y gnd NAND2X1_189/Y vdd NAND2X1
XNAND2X1_167 MUX2X1_1/B BUFX4_173/Y gnd AOI22X1_45/A vdd NAND2X1
XNAND2X1_123 MUX2X1_1/Y BUFX4_197/Y gnd AOI21X1_30/A vdd NAND2X1
XNAND2X1_156 INVX2_154/Y BUFX4_177/Y gnd AOI22X1_39/A vdd NAND2X1
XOAI21X1_651 OAI21X1_651/A OAI21X1_650/Y OAI21X1_651/C gnd DFFSR_148/D vdd OAI21X1
XOAI21X1_673 OAI21X1_673/A BUFX4_204/Y NAND2X1_294/Y gnd DFFSR_137/D vdd OAI21X1
XOAI21X1_640 NOR2X1_293/Y INVX2_76/Y BUFX4_120/Y gnd OAI21X1_640/Y vdd OAI21X1
XOAI21X1_684 BUFX4_58/Y NAND2X1_299/Y OAI21X1_684/C gnd OAI21X1_686/A vdd OAI21X1
XAOI21X1_4 AOI21X1_4/A AOI21X1_2/B AOI21X1_4/C gnd AOI21X1_4/Y vdd AOI21X1
XINVX2_4 INVX2_4/A gnd INVX2_4/Y vdd INVX2
XOAI21X1_662 NOR2X1_304/Y OAI21X1_662/B OAI21X1_662/C gnd DFFSR_141/D vdd OAI21X1
XXNOR2X1_12 OR2X2_8/A INVX4_11/A gnd XNOR2X1_12/Y vdd XNOR2X1
XOAI21X1_695 NOR2X1_315/Y OAI21X1_695/B OAI21X1_695/C gnd DFFSR_130/D vdd OAI21X1
XBUFX2_22 BUFX2_22/A gnd ss_pad_o[19] vdd BUFX2
XBUFX2_11 BUFX2_11/A gnd ss_pad_o[8] vdd BUFX2
XBUFX2_44 BUFX2_44/A gnd wb_dat_o[8] vdd BUFX2
XINVX1_80 DFFSR_98/Q gnd INVX1_80/Y vdd INVX1
XBUFX2_33 BUFX2_33/A gnd ss_pad_o[30] vdd BUFX2
XINVX1_91 INVX1_91/A gnd INVX1_91/Y vdd INVX1
XFILL_31_1_1 gnd vdd FILL
XBUFX2_55 BUFX2_55/A gnd wb_dat_o[19] vdd BUFX2
XBUFX2_66 BUFX2_66/A gnd wb_dat_o[30] vdd BUFX2
XNOR2X1_2 NOR2X1_2/A NOR2X1_2/B gnd NOR2X1_2/Y vdd NOR2X1
XAOI21X1_34 OR2X2_10/Y AOI21X1_34/B AOI21X1_33/Y gnd AOI21X1_34/Y vdd AOI21X1
XFILL_22_1_1 gnd vdd FILL
XAOI21X1_23 INVX2_41/Y AND2X2_8/A INVX1_75/Y gnd AOI21X1_23/Y vdd AOI21X1
XAOI21X1_12 INVX1_97/A BUFX4_190/Y AOI21X1_12/C gnd AOI21X1_12/Y vdd AOI21X1
XAOI21X1_45 AOI21X1_43/Y AOI21X1_45/B AND2X2_20/Y gnd AOI21X1_45/Y vdd AOI21X1
XAOI21X1_78 INVX2_94/Y BUFX4_174/Y INVX1_117/A gnd AOI22X1_51/C vdd AOI21X1
XAOI21X1_89 INVX2_117/Y BUFX4_174/Y INVX1_117/A gnd AOI21X1_89/Y vdd AOI21X1
XAOI21X1_67 AOI21X1_67/A AOI22X1_46/Y INVX1_125/A gnd NOR3X1_3/A vdd AOI21X1
XOAI21X1_7 INVX1_4/Y MUX2X1_7/S OAI21X1_7/C gnd NAND3X1_6/B vdd OAI21X1
XAOI21X1_56 INVX2_153/Y BUFX4_158/Y AOI21X1_69/C gnd AOI22X1_39/B vdd AOI21X1
XFILL_5_2_1 gnd vdd FILL
XOAI22X1_42 INVX2_46/Y BUFX4_101/Y OAI22X1_42/C OAI22X1_42/D gnd DFFSR_247/D vdd OAI22X1
XOAI22X1_20 OAI22X1_7/D INVX2_38/Y OAI22X1_4/C INVX1_45/Y gnd NOR2X1_11/B vdd OAI22X1
XOAI22X1_31 BUFX4_199/Y INVX2_27/Y OAI22X1_4/C INVX1_56/Y gnd NOR2X1_16/B vdd OAI22X1
XFILL_13_1_1 gnd vdd FILL
XOAI21X1_492 INVX2_101/Y BUFX4_160/Y NAND2X1_229/Y gnd OAI21X1_492/Y vdd OAI21X1
XOAI21X1_481 BUFX4_211/Y BUFX4_28/Y INVX2_79/A gnd OAI21X1_485/C vdd OAI21X1
XOAI21X1_470 BUFX4_220/Y OAI21X1_470/B BUFX4_48/Y gnd AOI21X1_164/A vdd OAI21X1
XBUFX4_139 INVX8_7/Y gnd DFFSR_1/R vdd BUFX4
XBUFX4_106 INVX8_4/Y gnd BUFX4_106/Y vdd BUFX4
XBUFX4_128 INVX8_24/Y gnd DFFSR_151/R vdd BUFX4
XBUFX4_117 INVX8_21/Y gnd BUFX4_117/Y vdd BUFX4
XFILL_1_1 gnd vdd FILL
XFILL_27_0_1 gnd vdd FILL
XFILL_2_0_1 gnd vdd FILL
XINVX2_106 DFFSR_180/Q gnd INVX2_106/Y vdd INVX2
XINVX2_117 AOI21X1_4/A gnd INVX2_117/Y vdd INVX2
XINVX2_128 INVX2_128/A gnd INVX2_128/Y vdd INVX2
XINVX2_139 DFFSR_141/Q gnd MUX2X1_2/B vdd INVX2
XFILL_18_0_1 gnd vdd FILL
XINVX1_161 INVX1_161/A gnd INVX1_161/Y vdd INVX1
XINVX1_150 INVX1_150/A gnd INVX1_150/Y vdd INVX1
XAOI21X1_121 INVX2_102/Y AOI21X1_121/B BUFX4_152/Y gnd OAI21X1_380/C vdd AOI21X1
XAOI21X1_110 NOR2X1_210/Y BUFX4_65/Y OAI21X1_352/Y gnd OAI21X1_355/A vdd AOI21X1
XAOI21X1_132 NOR2X1_222/Y BUFX4_67/Y AOI21X1_132/C gnd OAI21X1_400/A vdd AOI21X1
XAOI21X1_143 AOI21X1_142/Y OAI21X1_428/Y NOR2X1_229/Y gnd DFFSR_214/D vdd AOI21X1
XAOI21X1_187 NOR2X1_264/Y BUFX4_58/Y AOI21X1_187/C gnd AOI21X1_187/Y vdd AOI21X1
XAOI21X1_165 INVX2_91/Y OR2X2_15/Y INVX8_19/A gnd OAI21X1_472/C vdd AOI21X1
XAOI21X1_198 NOR2X1_272/Y BUFX4_63/Y AOI21X1_198/C gnd AOI21X1_198/Y vdd AOI21X1
XAOI21X1_154 NOR2X1_236/Y BUFX4_63/Y AOI21X1_154/C gnd OAI21X1_447/A vdd AOI21X1
XAOI21X1_176 INVX2_113/Y AOI21X1_176/B BUFX4_229/Y gnd OAI21X1_507/C vdd AOI21X1
XNAND3X1_114 INVX8_10/Y OAI21X1_210/Y OAI21X1_211/Y gnd NAND3X1_114/Y vdd NAND3X1
XNAND3X1_103 INVX1_66/Y INVX1_67/Y NOR2X1_32/Y gnd NOR2X1_34/A vdd NAND3X1
XNAND3X1_136 BUFX4_239/Y OAI21X1_234/Y NAND3X1_136/C gnd NAND3X1_137/C vdd NAND3X1
XNAND3X1_158 INVX4_4/A NAND3X1_158/B NAND3X1_157/Y gnd NAND3X1_159/C vdd NAND3X1
XNAND3X1_169 NOR2X1_51/Y NAND3X1_140/Y NAND3X1_169/C gnd NAND3X1_169/Y vdd NAND3X1
XNAND3X1_147 INVX2_47/A NAND3X1_143/Y NAND3X1_146/Y gnd NAND3X1_155/B vdd NAND3X1
XNAND3X1_125 BUFX4_195/Y NAND2X1_115/Y NAND2X1_116/Y gnd NAND3X1_125/Y vdd NAND3X1
XFILL_13_2 gnd vdd FILL
XDFFSR_134 INVX2_80/A CLKBUF1_12/A DFFSR_137/R vdd DFFSR_134/D gnd vdd DFFSR
XDFFSR_123 DFFSR_123/Q CLKBUF1_12/Y DFFSR_151/R vdd DFFSR_123/D gnd vdd DFFSR
XDFFSR_167 AOI22X1_7/A DFFSR_92/CLK DFFSR_167/R vdd DFFSR_167/D gnd vdd DFFSR
XDFFSR_156 INVX1_47/A CLKBUF1_50/Y DFFSR_167/R vdd DFFSR_156/D gnd vdd DFFSR
XBUFX4_8 wb_sel_i[1] gnd BUFX4_8/Y vdd BUFX4
XDFFSR_145 MUX2X1_5/B CLKBUF1_34/Y DFFSR_174/R vdd DFFSR_145/D gnd vdd DFFSR
XDFFSR_178 INVX2_64/A CLKBUF1_24/Y DFFSR_194/R vdd DFFSR_178/D gnd vdd DFFSR
XDFFSR_112 DFFSR_112/Q DFFSR_7/CLK vdd BUFX4_89/Y DFFSR_112/D gnd vdd DFFSR
XDFFSR_101 XOR2X1_1/B DFFSR_56/CLK vdd DFFSR_98/R DFFSR_101/D gnd vdd DFFSR
XDFFSR_189 DFFSR_189/Q CLKBUF1_39/Y DFFSR_203/R vdd DFFSR_189/D gnd vdd DFFSR
XNAND2X1_327 INVX8_23/A NOR2X1_312/Y gnd INVX1_161/A vdd NAND2X1
XNAND2X1_316 BUFX4_204/Y OAI21X1_715/Y gnd OAI21X1_717/C vdd NAND2X1
XNAND2X1_305 INVX8_22/A NOR2X1_312/Y gnd INVX1_153/A vdd NAND2X1
XNAND2X1_338 INVX8_22/A INVX1_164/A gnd NAND2X1_338/Y vdd NAND2X1
XINVX4_8 INVX4_8/A gnd INVX4_8/Y vdd INVX4
XFILL_35_6_0 gnd vdd FILL
XOAI21X1_129 BUFX4_93/Y BUFX4_103/Y DFFSR_3/Q gnd BUFX2_5/A vdd OAI21X1
XOAI21X1_118 INVX2_35/Y BUFX4_83/Y OAI21X1_86/C gnd NAND3X1_63/B vdd OAI21X1
XOAI21X1_107 AND2X2_3/Y INVX2_29/Y NAND3X1_57/Y gnd DFFSR_61/D vdd OAI21X1
XBUFX2_5 BUFX2_5/A gnd ss_pad_o[2] vdd BUFX2
XNAND2X1_102 INVX2_42/Y INVX1_86/A gnd OR2X2_7/A vdd NAND2X1
XNAND2X1_135 INVX4_2/Y NOR2X1_175/B gnd NAND2X1_136/B vdd NAND2X1
XNAND2X1_146 NAND2X1_145/Y NOR2X1_179/Y gnd AOI21X1_54/C vdd NAND2X1
XNAND2X1_113 INVX2_54/Y NOR2X1_97/B gnd NAND3X1_109/C vdd NAND2X1
XNAND2X1_179 INVX2_95/Y BUFX4_156/Y gnd AOI22X1_51/D vdd NAND2X1
XNAND2X1_168 MUX2X1_4/B BUFX4_153/Y gnd AOI22X1_45/D vdd NAND2X1
XNAND2X1_124 MUX2X1_2/Y BUFX4_188/Y gnd AOI21X1_30/B vdd NAND2X1
XNAND2X1_157 INVX2_155/Y BUFX4_158/Y gnd AOI22X1_39/D vdd NAND2X1
XFILL_26_6_0 gnd vdd FILL
XNOR2X1_190 INVX1_114/A INVX1_113/Y gnd NOR2X1_190/Y vdd NOR2X1
XFILL_1_6_0 gnd vdd FILL
XOAI21X1_641 INVX2_76/Y BUFX4_80/Y NAND2X1_244/Y gnd OAI21X1_641/Y vdd OAI21X1
XOAI21X1_685 INVX2_80/Y BUFX4_165/Y NAND2X1_224/Y gnd OAI21X1_685/Y vdd OAI21X1
XAOI21X1_5 INVX2_94/A AOI21X1_7/B AOI21X1_5/C gnd AOI21X1_5/Y vdd AOI21X1
XOAI21X1_630 BUFX4_58/Y OR2X2_17/Y AOI21X1_230/Y gnd AOI21X1_232/B vdd OAI21X1
XOAI21X1_674 INVX2_90/Y BUFX4_163/Y NAND2X1_219/Y gnd NAND2X1_295/B vdd OAI21X1
XINVX2_5 INVX2_5/A gnd INVX2_5/Y vdd INVX2
XOAI21X1_652 INVX1_92/Y BUFX4_72/Y OAI21X1_323/C gnd NAND2X1_283/B vdd OAI21X1
XOAI21X1_663 INVX1_120/Y BUFX4_71/Y OAI21X1_353/C gnd NAND2X1_289/B vdd OAI21X1
XOAI21X1_696 INVX2_156/Y BUFX4_8/Y NAND2X1_232/Y gnd NAND2X1_307/B vdd OAI21X1
XBUFX2_56 DFFSR_85/Q gnd wb_dat_o[20] vdd BUFX2
XBUFX2_23 BUFX2_23/A gnd ss_pad_o[20] vdd BUFX2
XINVX1_81 INVX1_81/A gnd INVX1_81/Y vdd INVX1
XBUFX2_45 DFFSR_74/Q gnd wb_dat_o[9] vdd BUFX2
XBUFX2_12 BUFX2_12/A gnd ss_pad_o[9] vdd BUFX2
XFILL_17_6_0 gnd vdd FILL
XINVX1_92 INVX1_92/A gnd INVX1_92/Y vdd INVX1
XBUFX2_67 BUFX2_67/A gnd wb_dat_o[31] vdd BUFX2
XBUFX2_34 BUFX2_34/A gnd ss_pad_o[31] vdd BUFX2
XINVX1_70 INVX1_70/A gnd INVX1_70/Y vdd INVX1
XNOR2X1_3 wb_adr_i[2] wb_adr_i[3] gnd NOR2X1_3/Y vdd NOR2X1
XAOI21X1_46 AOI21X1_46/A OR2X2_7/A INVX8_13/A gnd AOI21X1_46/Y vdd AOI21X1
XAOI21X1_35 INVX4_3/A AOI21X1_35/B AOI21X1_43/B gnd AOI21X1_35/Y vdd AOI21X1
XAOI21X1_13 INVX2_87/A AOI21X1_7/B AOI21X1_13/C gnd NAND2X1_56/A vdd AOI21X1
XAOI21X1_68 INVX1_119/Y OR2X2_3/B AOI21X1_68/C gnd NOR3X1_3/B vdd AOI21X1
XAOI21X1_24 OR2X2_5/B OR2X2_5/A BUFX4_2/Y gnd AOI21X1_24/Y vdd AOI21X1
XAOI21X1_57 INVX2_156/Y BUFX4_177/Y INVX1_117/A gnd AOI22X1_39/C vdd AOI21X1
XAOI21X1_79 INVX2_89/Y BUFX4_155/Y AOI21X1_71/C gnd AOI21X1_79/Y vdd AOI21X1
XOAI21X1_8 BUFX4_180/Y INVX1_4/Y OAI21X1_8/C gnd DFFSR_28/D vdd OAI21X1
XOAI22X1_43 INVX4_2/Y BUFX4_101/Y OAI22X1_43/C OAI22X1_43/D gnd DFFSR_248/D vdd OAI22X1
XOAI22X1_10 INVX8_1/A INVX2_13/Y INVX2_35/Y OAI22X1_7/D gnd NOR2X1_8/A vdd OAI22X1
XOAI22X1_21 BUFX4_76/Y INVX2_1/Y INVX1_46/Y INVX8_6/A gnd NOR2X1_12/A vdd OAI22X1
XOAI22X1_32 BUFX4_76/Y INVX2_6/Y INVX2_28/Y INVX8_4/A gnd NOR2X1_17/A vdd OAI22X1
XOAI21X1_493 BUFX4_220/Y OAI21X1_492/Y BUFX4_47/Y gnd AOI21X1_171/A vdd OAI21X1
XOAI21X1_482 NOR2X1_250/Y INVX2_79/Y BUFX4_170/Y gnd OAI21X1_482/Y vdd OAI21X1
XOAI21X1_471 BUFX4_98/Y INVX4_6/Y INVX1_127/Y gnd OR2X2_15/A vdd OAI21X1
XOAI21X1_460 BUFX4_205/Y BUFX4_29/Y DFFSR_204/Q gnd OAI21X1_460/Y vdd OAI21X1
XFILL_32_4_0 gnd vdd FILL
XFILL_23_4_0 gnd vdd FILL
XBUFX4_107 INVX8_4/Y gnd BUFX4_107/Y vdd BUFX4
XFILL_6_5_0 gnd vdd FILL
XBUFX4_118 INVX8_21/Y gnd BUFX4_118/Y vdd BUFX4
XBUFX4_129 INVX8_24/Y gnd DFFSR_203/R vdd BUFX4
XFILL_14_4_0 gnd vdd FILL
XOAI21X1_290 AOI21X1_45/Y NOR2X1_178/Y NOR2X1_179/Y gnd AOI21X1_53/B vdd OAI21X1
XFILL_1_2 gnd vdd FILL
XFILL_36_1 gnd vdd FILL
XINVX2_107 DFFSR_116/Q gnd INVX2_107/Y vdd INVX2
XINVX2_118 DFFSR_199/Q gnd INVX2_118/Y vdd INVX2
XINVX2_129 INVX2_129/A gnd INVX2_129/Y vdd INVX2
XDFFSR_90 BUFX2_61/A CLKBUF1_34/A DFFSR_25/R vdd DFFSR_90/D gnd vdd DFFSR
XINVX1_151 INVX1_151/A gnd INVX1_151/Y vdd INVX1
XINVX1_162 INVX1_162/A gnd INVX1_162/Y vdd INVX1
XINVX1_140 INVX1_140/A gnd INVX1_140/Y vdd INVX1
XAOI21X1_122 BUFX4_151/Y OAI21X1_381/Y BUFX4_47/Y gnd AOI21X1_123/A vdd AOI21X1
XAOI21X1_100 INVX2_56/Y BUFX4_176/Y INVX1_118/A gnd AOI21X1_100/Y vdd AOI21X1
XAOI21X1_144 INVX2_145/Y OR2X2_13/Y BUFX4_152/Y gnd AOI21X1_144/Y vdd AOI21X1
XAOI21X1_111 NOR2X1_211/Y BUFX4_66/Y AOI21X1_111/C gnd OAI21X1_360/A vdd AOI21X1
XFILL_20_2_0 gnd vdd FILL
XAOI21X1_166 AOI21X1_166/A AOI21X1_166/B NOR2X1_247/Y gnd DFFSR_200/D vdd AOI21X1
XAOI21X1_155 INVX2_110/Y NAND2X1_249/Y BUFX4_231/Y gnd OAI21X1_449/C vdd AOI21X1
XAOI21X1_133 NOR2X1_223/Y BUFX4_67/Y AOI21X1_133/C gnd OAI21X1_405/A vdd AOI21X1
XAOI21X1_188 AND2X2_27/Y BUFX4_61/Y OAI21X1_554/Y gnd AOI21X1_188/Y vdd AOI21X1
XAOI21X1_199 NOR2X1_273/Y BUFX4_57/Y OAI21X1_581/Y gnd OAI21X1_584/A vdd AOI21X1
XAOI21X1_177 AOI21X1_177/A AOI21X1_177/B NOR2X1_258/Y gnd DFFSR_191/D vdd AOI21X1
XFILL_28_3_0 gnd vdd FILL
XNAND3X1_137 INVX4_4/A NAND3X1_135/Y NAND3X1_137/C gnd NAND3X1_138/C vdd NAND3X1
XFILL_3_3_0 gnd vdd FILL
XNAND3X1_126 INVX8_10/Y NAND3X1_125/Y OAI21X1_220/Y gnd NAND3X1_128/B vdd NAND3X1
XNAND3X1_148 MUX2X1_1/S NAND3X1_148/B OAI21X1_245/Y gnd NAND3X1_148/Y vdd NAND3X1
XNAND3X1_115 INVX4_4/Y NAND3X1_113/Y NAND3X1_114/Y gnd NAND3X1_115/Y vdd NAND3X1
XNAND3X1_104 INVX1_68/Y INVX1_69/Y NOR2X1_33/Y gnd NOR2X1_34/B vdd NAND3X1
XNAND3X1_159 INVX2_47/A OAI21X1_252/Y NAND3X1_159/C gnd NAND3X1_159/Y vdd NAND3X1
XFILL_11_2_0 gnd vdd FILL
XFILL_19_3_0 gnd vdd FILL
XDFFSR_168 INVX2_88/A DFFSR_78/CLK DFFSR_151/R vdd DFFSR_168/D gnd vdd DFFSR
XDFFSR_135 DFFSR_135/Q CLKBUF1_5/A DFFSR_130/R vdd DFFSR_135/D gnd vdd DFFSR
XBUFX4_9 wb_sel_i[1] gnd BUFX4_9/Y vdd BUFX4
XDFFSR_146 INVX1_92/A DFFSR_26/CLK DFFSR_174/R vdd DFFSR_146/D gnd vdd DFFSR
XDFFSR_179 INVX2_126/A CLKBUF1_34/A DFFSR_174/R vdd DFFSR_179/D gnd vdd DFFSR
XDFFSR_113 OR2X2_6/B DFFSR_98/CLK vdd BUFX4_87/Y DFFSR_113/D gnd vdd DFFSR
XDFFSR_124 INVX2_96/A CLKBUF1_8/Y DFFSR_130/R vdd DFFSR_124/D gnd vdd DFFSR
XDFFSR_102 INVX1_70/A DFFSR_87/CLK vdd DFFSR_98/R DFFSR_102/D gnd vdd DFFSR
XDFFSR_157 INVX1_49/A CLKBUF1_45/Y DFFSR_167/R vdd DFFSR_157/D gnd vdd DFFSR
XNAND2X1_317 INVX8_23/A NOR2X1_308/Y gnd INVX1_158/A vdd NAND2X1
XNAND2X1_339 BUFX4_206/Y NAND2X1_339/B gnd OAI21X1_786/C vdd NAND2X1
XNAND2X1_306 BUFX4_205/Y NAND2X1_306/B gnd OAI21X1_695/C vdd NAND2X1
XNAND2X1_328 BUFX4_6/Y wb_dat_i[15] gnd NAND2X1_328/Y vdd NAND2X1
XNOR2X1_350 INVX4_5/A DFFSR_41/Q gnd NOR2X1_350/Y vdd NOR2X1
XINVX4_9 INVX4_9/A gnd INVX4_9/Y vdd INVX4
XFILL_35_6_1 gnd vdd FILL
XFILL_34_1_0 gnd vdd FILL
XNAND3X1_90 NAND2X1_64/Y AOI22X1_9/Y NAND3X1_90/C gnd DFFSR_85/D vdd NAND3X1
XNOR2X1_90 INVX1_94/Y BUFX4_40/Y gnd NOR2X1_90/Y vdd NOR2X1
XOAI21X1_119 AND2X2_3/Y INVX2_35/Y NAND3X1_63/Y gnd DFFSR_51/D vdd OAI21X1
XOAI21X1_108 INVX2_30/Y BUFX4_10/Y OAI21X1_47/C gnd NAND3X1_58/B vdd OAI21X1
XNAND2X1_114 INVX8_9/Y INVX1_90/Y gnd OAI21X1_204/C vdd NAND2X1
XBUFX2_6 BUFX2_6/A gnd ss_pad_o[3] vdd BUFX2
XNAND2X1_103 DFFSR_43/Q INVX1_80/Y gnd NAND2X1_103/Y vdd NAND2X1
XNAND2X1_125 MUX2X1_3/Y AND2X2_16/B gnd AOI21X1_31/A vdd NAND2X1
XNAND2X1_136 NAND2X1_136/A NAND2X1_136/B gnd OAI21X1_273/B vdd NAND2X1
XNAND2X1_147 OR2X2_8/B INVX8_13/Y gnd AOI21X1_44/A vdd NAND2X1
XNAND2X1_1 wb_dat_i[24] MUX2X1_7/S gnd OAI21X1_1/C vdd NAND2X1
XNAND2X1_158 INVX2_151/Y BUFX4_177/Y gnd AOI22X1_40/A vdd NAND2X1
XNAND2X1_169 AOI22X1_44/Y AOI22X1_45/Y gnd AOI22X1_46/D vdd NAND2X1
XNOR2X1_180 INVX4_3/Y NOR2X1_180/B gnd NOR2X1_180/Y vdd NOR2X1
XFILL_26_6_1 gnd vdd FILL
XFILL_25_1_0 gnd vdd FILL
XINVX2_6 INVX2_6/A gnd INVX2_6/Y vdd INVX2
XNOR2X1_191 INVX1_114/Y INVX1_113/A gnd NOR2X1_191/Y vdd NOR2X1
XFILL_1_6_1 gnd vdd FILL
XFILL_0_1_0 gnd vdd FILL
XAOI21X1_6 DFFSR_121/Q AOI21X1_2/B AOI21X1_6/C gnd AOI21X1_6/Y vdd AOI21X1
XOAI21X1_642 BUFX4_120/Y OAI21X1_641/Y BUFX4_114/Y gnd OAI21X1_642/Y vdd OAI21X1
XOAI21X1_686 OAI21X1_686/A BUFX4_206/Y NAND2X1_301/Y gnd DFFSR_134/D vdd OAI21X1
XOAI21X1_631 INVX2_58/Y BUFX4_84/Y NAND2X1_239/Y gnd AOI21X1_231/B vdd OAI21X1
XOAI21X1_675 BUFX4_98/Y INVX8_18/Y NOR2X1_276/Y gnd INVX1_150/A vdd OAI21X1
XOAI21X1_653 BUFX4_96/Y INVX8_18/Y AND2X2_28/A gnd NOR2X1_296/B vdd OAI21X1
XOAI21X1_664 NOR2X1_1/A INVX8_18/Y INVX1_140/Y gnd OR2X2_19/A vdd OAI21X1
XOAI21X1_620 BUFX4_57/Y AOI21X1_220/B OAI21X1_620/C gnd AOI21X1_222/B vdd OAI21X1
XOAI21X1_697 INVX1_155/A DFFSR_129/Q BUFX4_118/Y gnd OAI21X1_698/B vdd OAI21X1
XFILL_8_2_0 gnd vdd FILL
XINVX1_60 INVX2_63/A gnd INVX1_60/Y vdd INVX1
XBUFX2_57 DFFSR_86/Q gnd wb_dat_o[21] vdd BUFX2
XBUFX2_24 BUFX2_24/A gnd ss_pad_o[21] vdd BUFX2
XBUFX2_35 BUFX2_35/A gnd wb_ack_o vdd BUFX2
XINVX1_82 INVX1_82/A gnd INVX1_82/Y vdd INVX1
XFILL_17_6_1 gnd vdd FILL
XFILL_16_1_0 gnd vdd FILL
XBUFX2_68 gnd gnd wb_err_o vdd BUFX2
XINVX1_71 DFFSR_51/Q gnd INVX1_71/Y vdd INVX1
XINVX1_93 INVX1_93/A gnd INVX1_93/Y vdd INVX1
XBUFX2_13 BUFX2_13/A gnd ss_pad_o[10] vdd BUFX2
XBUFX2_46 BUFX2_46/A gnd wb_dat_o[10] vdd BUFX2
XNOR2X1_4 wb_adr_i[4] wb_adr_i[2] gnd NOR2X1_4/Y vdd NOR2X1
XAOI21X1_36 INVX8_13/A AOI21X1_36/B INVX2_42/Y gnd AOI21X1_36/Y vdd AOI21X1
XAOI21X1_47 INVX2_48/A BUFX4_112/Y INVX2_18/A gnd AOI21X1_47/Y vdd AOI21X1
XAOI21X1_69 INVX2_104/Y BUFX4_154/Y AOI21X1_69/C gnd AOI21X1_69/Y vdd AOI21X1
XAOI21X1_58 INVX2_150/Y BUFX4_158/Y AOI21X1_71/C gnd AOI21X1_58/Y vdd AOI21X1
XAOI21X1_25 OR2X2_6/B OR2X2_6/A BUFX4_4/Y gnd AOI22X1_35/D vdd AOI21X1
XAOI21X1_14 DFFSR_129/Q BUFX4_190/Y OAI22X1_34/Y gnd NAND2X1_57/A vdd AOI21X1
XOAI21X1_9 INVX1_5/Y BUFX4_70/Y OAI21X1_9/C gnd NAND3X1_7/B vdd OAI21X1
XOAI22X1_44 INVX4_3/Y BUFX4_101/Y OAI22X1_44/C NOR2X1_342/Y gnd DFFSR_249/D vdd OAI22X1
XOAI22X1_11 OAI22X1_4/C INVX1_35/Y INVX1_36/Y INVX8_5/A gnd NOR2X1_8/B vdd OAI22X1
XOAI22X1_22 INVX8_4/A INVX2_23/Y OAI22X1_4/C INVX1_47/Y gnd NOR2X1_12/B vdd OAI22X1
XOAI21X1_450 INVX2_110/Y MUX2X1_7/S OAI21X1_567/C gnd OAI21X1_451/B vdd OAI21X1
XOAI22X1_33 OAI22X1_4/C INVX1_57/Y INVX1_58/Y INVX8_5/A gnd NOR2X1_17/B vdd OAI22X1
XOAI21X1_483 INVX2_79/Y BUFX4_165/Y NAND2X1_224/Y gnd OAI21X1_484/B vdd OAI21X1
XOAI21X1_472 BUFX4_59/Y OR2X2_15/Y OAI21X1_472/C gnd AOI21X1_166/B vdd OAI21X1
XOAI21X1_494 BUFX4_67/Y AOI21X1_172/B OAI21X1_494/C gnd AOI21X1_173/B vdd OAI21X1
XOAI21X1_461 NOR2X1_242/Y INVX1_135/Y BUFX4_167/Y gnd AOI21X1_160/C vdd OAI21X1
XFILL_32_4_1 gnd vdd FILL
XFILL_23_4_1 gnd vdd FILL
XBUFX4_108 INVX8_4/Y gnd BUFX4_108/Y vdd BUFX4
XFILL_5_0_0 gnd vdd FILL
XFILL_6_5_1 gnd vdd FILL
XBUFX4_119 INVX8_20/Y gnd BUFX4_119/Y vdd BUFX4
XFILL_14_4_1 gnd vdd FILL
XOAI21X1_280 INVX1_107/Y BUFX4_112/Y AOI21X1_47/Y gnd NAND2X1_150/A vdd OAI21X1
XOAI21X1_291 AOI21X1_53/Y INVX1_106/A AND2X2_21/Y gnd INVX1_117/A vdd OAI21X1
XFILL_36_2 gnd vdd FILL
XFILL_29_1 gnd vdd FILL
XINVX2_119 DFFSR_135/Q gnd INVX2_119/Y vdd INVX2
XINVX2_108 DFFSR_239/Q gnd INVX2_108/Y vdd INVX2
XDFFSR_91 BUFX2_62/A DFFSR_61/CLK DFFSR_95/R vdd DFFSR_91/D gnd vdd DFFSR
XDFFSR_80 BUFX2_51/A CLKBUF1_2/Y DFFSR_25/R vdd DFFSR_80/D gnd vdd DFFSR
XINVX1_152 INVX1_152/A gnd INVX1_152/Y vdd INVX1
XINVX1_141 INVX1_141/A gnd INVX1_141/Y vdd INVX1
XINVX1_130 INVX1_130/A gnd INVX1_130/Y vdd INVX1
XINVX1_163 INVX1_163/A gnd INVX1_163/Y vdd INVX1
XAOI21X1_123 AOI21X1_123/A OAI21X1_380/Y NOR2X1_217/Y gnd DFFSR_228/D vdd AOI21X1
XAOI21X1_145 BUFX4_151/Y OAI21X1_431/Y BUFX4_47/Y gnd AOI21X1_146/A vdd AOI21X1
XAOI21X1_101 INVX2_60/Y BUFX4_176/Y INVX1_117/A gnd AOI21X1_101/Y vdd AOI21X1
XFILL_20_2_1 gnd vdd FILL
XAOI21X1_167 NOR2X1_248/Y BUFX4_60/Y AOI21X1_167/C gnd OAI21X1_480/A vdd AOI21X1
XAOI21X1_112 NOR2X1_212/Y BUFX4_59/Y OAI21X1_362/Y gnd OAI21X1_365/A vdd AOI21X1
XAOI21X1_189 AND2X2_28/Y BUFX4_65/Y OAI21X1_558/Y gnd OAI21X1_561/A vdd AOI21X1
XAOI21X1_156 AOI21X1_156/A AOI21X1_156/B NOR2X1_237/Y gnd DFFSR_207/D vdd AOI21X1
XAOI21X1_178 INVX2_72/Y NAND2X1_256/Y BUFX4_229/Y gnd OAI21X1_510/C vdd AOI21X1
XAOI21X1_134 NOR2X1_224/Y BUFX4_67/Y AOI21X1_134/C gnd OAI21X1_410/A vdd AOI21X1
XFILL_28_3_1 gnd vdd FILL
XFILL_3_3_1 gnd vdd FILL
XNAND3X1_138 INVX2_47/A NAND3X1_133/Y NAND3X1_138/C gnd NAND3X1_139/B vdd NAND3X1
XNAND3X1_116 INVX2_47/Y NAND3X1_116/B NAND3X1_115/Y gnd NAND3X1_124/B vdd NAND3X1
XNAND3X1_105 NOR2X1_35/Y NOR2X1_36/Y NOR2X1_37/Y gnd NOR2X1_38/B vdd NAND3X1
XNAND3X1_127 BUFX4_237/Y OAI21X1_221/Y OAI21X1_222/Y gnd NAND3X1_128/C vdd NAND3X1
XNAND3X1_149 INVX8_10/Y OAI21X1_246/Y OAI21X1_247/Y gnd NAND3X1_149/Y vdd NAND3X1
XFILL_11_2_1 gnd vdd FILL
XFILL_19_3_1 gnd vdd FILL
XDFFSR_114 DFFSR_114/Q DFFSR_99/CLK vdd BUFX4_87/Y DFFSR_114/D gnd vdd DFFSR
XDFFSR_103 DFFSR_103/Q DFFSR_28/CLK vdd BUFX4_90/Y DFFSR_103/D gnd vdd DFFSR
XDFFSR_125 INVX2_138/A CLKBUF1_1/Y DFFSR_130/R vdd DFFSR_125/D gnd vdd DFFSR
XDFFSR_169 DFFSR_169/Q CLKBUF1_5/Y DFFSR_137/R vdd DFFSR_169/D gnd vdd DFFSR
XNAND2X1_318 BUFX4_208/Y OAI21X1_718/Y gnd NAND2X1_318/Y vdd NAND2X1
XDFFSR_136 INVX2_90/A CLKBUF1_19/Y DFFSR_151/R vdd DFFSR_136/D gnd vdd DFFSR
XDFFSR_147 AND2X2_17/B CLKBUF1_28/Y DFFSR_174/R vdd DFFSR_147/D gnd vdd DFFSR
XDFFSR_158 INVX1_51/A DFFSR_98/CLK DFFSR_130/R vdd DFFSR_158/D gnd vdd DFFSR
XNAND2X1_307 BUFX4_210/Y NAND2X1_307/B gnd NAND2X1_307/Y vdd NAND2X1
XNAND2X1_329 INVX1_111/A NOR2X1_190/Y gnd OR2X2_21/B vdd NAND2X1
XNOR2X1_340 INVX4_11/Y INVX2_45/Y gnd OAI22X1_42/C vdd NOR2X1
XNAND3X1_91 AOI22X1_12/Y NAND3X1_91/B AOI22X1_11/Y gnd DFFSR_86/D vdd NAND3X1
XNAND3X1_80 wb_adr_i[3] DFFSR_189/Q NOR2X1_4/Y gnd NAND3X1_80/Y vdd NAND3X1
XFILL_34_1_1 gnd vdd FILL
XNOR2X1_91 INVX2_73/Y BUFX4_217/Y gnd NOR2X1_91/Y vdd NOR2X1
XNOR2X1_80 INVX2_65/Y NOR2X1_99/B gnd NOR2X1_80/Y vdd NOR2X1
XBUFX2_7 BUFX2_7/A gnd ss_pad_o[4] vdd BUFX2
XOAI21X1_109 AND2X2_3/Y INVX2_30/Y NAND3X1_58/Y gnd DFFSR_62/D vdd OAI21X1
XNAND2X1_137 OAI21X1_272/Y NOR2X1_177/B gnd AOI21X1_35/B vdd NAND2X1
XNAND2X1_104 OAI21X1_187/Y NOR2X1_48/B gnd NAND2X1_104/Y vdd NAND2X1
XNAND2X1_148 NAND2X1_148/A NAND2X1_148/B gnd INVX1_108/A vdd NAND2X1
XNAND2X1_159 INVX2_152/Y BUFX4_158/Y gnd AOI22X1_40/D vdd NAND2X1
XNAND2X1_115 INVX2_81/Y BUFX4_40/Y gnd NAND2X1_115/Y vdd NAND2X1
XNAND2X1_126 MUX2X1_4/Y AND2X2_15/B gnd AOI21X1_31/B vdd NAND2X1
XFILL_25_1_1 gnd vdd FILL
XNAND2X1_2 BUFX4_70/Y wb_dat_i[25] gnd OAI21X1_3/C vdd NAND2X1
XOAI21X1_610 BUFX4_122/Y OAI21X1_609/Y BUFX4_113/Y gnd OAI21X1_610/Y vdd OAI21X1
XNOR2X1_181 DFFSR_33/Q OR2X2_10/A gnd NOR2X1_181/Y vdd NOR2X1
XOAI21X1_632 NOR2X1_290/Y INVX2_159/Y BUFX4_121/Y gnd AOI21X1_233/C vdd OAI21X1
XINVX2_7 INVX2_7/A gnd INVX2_7/Y vdd INVX2
XNOR2X1_170 INVX2_160/Y NOR2X1_71/B gnd NOR2X1_170/Y vdd NOR2X1
XNOR2X1_192 BUFX4_156/Y INVX1_118/A gnd INVX8_22/A vdd NOR2X1
XFILL_0_1_1 gnd vdd FILL
XOAI21X1_621 INVX2_112/Y BUFX4_11/Y OAI21X1_621/C gnd AOI21X1_221/B vdd OAI21X1
XOAI21X1_687 INVX1_100/Y NAND2X1_9/B NAND2X1_226/Y gnd NAND2X1_302/B vdd OAI21X1
XOAI21X1_643 OAI21X1_643/A OAI21X1_642/Y NAND2X1_280/Y gnd DFFSR_150/D vdd OAI21X1
XAOI21X1_7 INVX2_60/A AOI21X1_7/B AOI21X1_7/C gnd AOI21X1_7/Y vdd AOI21X1
XOAI21X1_676 INVX1_150/A INVX8_22/Y INVX2_90/Y gnd OAI21X1_677/C vdd OAI21X1
XOAI21X1_665 INVX1_148/A INVX1_120/A BUFX4_117/Y gnd OAI21X1_665/Y vdd OAI21X1
XOAI21X1_654 INVX1_141/A INVX1_92/A BUFX4_117/Y gnd OAI21X1_655/B vdd OAI21X1
XOAI21X1_698 NOR2X1_317/Y OAI21X1_698/B NAND2X1_307/Y gnd DFFSR_129/D vdd OAI21X1
XINVX1_83 INVX1_83/A gnd INVX1_83/Y vdd INVX1
XINVX1_72 INVX1_72/A gnd INVX1_72/Y vdd INVX1
XFILL_8_2_1 gnd vdd FILL
XINVX1_94 INVX1_94/A gnd INVX1_94/Y vdd INVX1
XINVX1_50 INVX1_50/A gnd INVX1_50/Y vdd INVX1
XINVX1_61 INVX1_61/A gnd INVX1_61/Y vdd INVX1
XBUFX2_36 DFFSR_65/Q gnd wb_dat_o[0] vdd BUFX2
XBUFX2_69 DFFSR_63/Q gnd wb_int_o vdd BUFX2
XBUFX2_25 BUFX2_25/A gnd ss_pad_o[22] vdd BUFX2
XBUFX2_58 BUFX2_58/A gnd wb_dat_o[22] vdd BUFX2
XBUFX2_14 BUFX2_14/A gnd ss_pad_o[11] vdd BUFX2
XBUFX2_47 BUFX2_47/A gnd wb_dat_o[11] vdd BUFX2
XFILL_16_1_1 gnd vdd FILL
XNOR2X1_5 NOR2X1_5/A NOR2X1_5/B gnd NOR2X1_5/Y vdd NOR2X1
XAOI21X1_37 AND2X2_20/A AND2X2_20/B AOI21X1_37/C gnd AOI21X1_37/Y vdd AOI21X1
XAOI21X1_48 INVX1_108/Y AOI21X1_48/B INVX8_9/Y gnd AOI21X1_48/Y vdd AOI21X1
XAOI21X1_59 INVX1_101/Y BUFX4_177/Y INVX1_118/A gnd AOI22X1_40/C vdd AOI21X1
XAOI21X1_26 INVX1_78/A NOR2X1_44/Y BUFX4_4/Y gnd AOI21X1_27/B vdd AOI21X1
XAOI21X1_15 INVX2_61/A BUFX4_127/Y AOI21X1_15/C gnd NAND2X1_58/B vdd AOI21X1
XOAI22X1_12 OAI22X1_1/D INVX1_37/Y INVX8_2/A INVX2_20/Y gnd AOI21X1_5/C vdd OAI22X1
XOAI22X1_23 BUFX4_77/Y INVX2_2/Y INVX1_48/Y INVX8_6/A gnd NOR2X1_13/A vdd OAI22X1
XOAI22X1_34 BUFX4_226/Y INVX1_59/Y INVX8_2/A BUFX4_94/Y gnd OAI22X1_34/Y vdd OAI22X1
XOAI22X1_45 INVX2_50/Y BUFX4_101/Y OAI22X1_45/C OAI22X1_45/D gnd DFFSR_251/D vdd OAI22X1
XOAI21X1_484 BUFX4_170/Y OAI21X1_484/B BUFX4_36/Y gnd OAI21X1_485/B vdd OAI21X1
XOAI21X1_473 INVX2_91/Y BUFX4_163/Y NAND2X1_219/Y gnd OAI21X1_474/B vdd OAI21X1
XOAI21X1_440 INVX2_152/Y BUFX4_73/Y OAI21X1_328/C gnd OAI21X1_440/Y vdd OAI21X1
XOAI21X1_451 BUFX4_224/Y OAI21X1_451/B BUFX4_50/Y gnd AOI21X1_156/A vdd OAI21X1
XOAI21X1_462 INVX1_135/Y BUFX4_71/Y OAI21X1_353/C gnd OAI21X1_462/Y vdd OAI21X1
XOAI21X1_495 INVX2_63/Y BUFX4_9/Y NAND2X1_231/Y gnd OAI21X1_496/B vdd OAI21X1
XBUFX4_109 DFFSR_42/Q gnd INVX1_17/A vdd BUFX4
XFILL_5_0_1 gnd vdd FILL
XOAI21X1_270 NOR2X1_176/A INVX8_13/Y INVX2_43/A gnd OAI21X1_271/C vdd OAI21X1
XOAI21X1_292 AOI21X1_54/Y INVX1_116/Y INVX1_105/Y gnd NAND3X1_198/C vdd OAI21X1
XOAI21X1_281 OAI21X1_273/B AOI21X1_34/Y NAND2X1_136/A gnd AOI21X1_48/B vdd OAI21X1
XFILL_36_3 gnd vdd FILL
XINVX2_109 INVX2_109/A gnd INVX2_109/Y vdd INVX2
XDFFSR_70 DFFSR_70/Q DFFSR_85/CLK DFFSR_88/R vdd DFFSR_70/D gnd vdd DFFSR
XDFFSR_81 DFFSR_81/Q DFFSR_6/CLK DFFSR_88/R vdd DFFSR_81/D gnd vdd DFFSR
XDFFSR_92 DFFSR_92/Q DFFSR_92/CLK DFFSR_25/R vdd DFFSR_92/D gnd vdd DFFSR
XINVX1_153 INVX1_153/A gnd INVX1_153/Y vdd INVX1
XINVX1_164 INVX1_164/A gnd INVX1_164/Y vdd INVX1
XINVX1_142 INVX1_142/A gnd INVX1_142/Y vdd INVX1
XINVX1_120 INVX1_120/A gnd INVX1_120/Y vdd INVX1
XINVX1_131 INVX1_131/A gnd INVX1_131/Y vdd INVX1
XAOI21X1_168 NOR2X1_250/Y BUFX4_66/Y OAI21X1_482/Y gnd AOI21X1_168/Y vdd AOI21X1
XAOI21X1_146 AOI21X1_146/A AOI21X1_146/B NOR2X1_230/Y gnd DFFSR_213/D vdd AOI21X1
XAOI21X1_113 INVX2_89/Y NAND2X1_218/Y INVX8_15/A gnd OAI21X1_366/C vdd AOI21X1
XAOI21X1_135 NOR2X1_225/Y BUFX4_59/Y AOI21X1_135/C gnd OAI21X1_415/A vdd AOI21X1
XAOI21X1_157 AND2X2_23/Y BUFX4_63/Y AOI21X1_157/C gnd OAI21X1_456/A vdd AOI21X1
XAOI21X1_179 AOI21X1_179/A AOI21X1_179/B NOR2X1_259/Y gnd DFFSR_190/D vdd AOI21X1
XAOI21X1_124 INVX2_62/Y NAND2X1_230/Y BUFX4_148/Y gnd AOI21X1_124/Y vdd AOI21X1
XAOI21X1_102 AOI22X1_77/Y NOR3X1_3/Y NOR2X1_200/Y gnd BUFX4_61/A vdd AOI21X1
XNAND3X1_139 INVX1_84/A NAND3X1_139/B NAND3X1_139/C gnd NAND3X1_140/B vdd NAND3X1
XNAND3X1_128 INVX4_4/Y NAND3X1_128/B NAND3X1_128/C gnd NAND3X1_128/Y vdd NAND3X1
XNAND3X1_117 INVX8_10/Y OAI21X1_212/Y NAND3X1_117/C gnd NAND3X1_117/Y vdd NAND3X1
XNAND3X1_106 NOR2X1_1/A NOR2X1_40/Y NOR2X1_27/Y gnd NAND2X1_85/B vdd NAND3X1
XDFFSR_148 INVX1_27/A DFFSR_88/CLK DFFSR_165/R vdd DFFSR_148/D gnd vdd DFFSR
XDFFSR_137 DFFSR_137/Q DFFSR_2/CLK DFFSR_137/R vdd DFFSR_137/D gnd vdd DFFSR
XFILL_30_5_0 gnd vdd FILL
XDFFSR_104 INVX1_72/A CLKBUF1_8/A vdd BUFX4_89/Y DFFSR_104/D gnd vdd DFFSR
XDFFSR_126 INVX1_94/A CLKBUF1_52/Y DFFSR_130/R vdd DFFSR_126/D gnd vdd DFFSR
XDFFSR_115 INVX1_77/A CLKBUF1_35/Y vdd BUFX4_90/Y DFFSR_115/D gnd vdd DFFSR
XNAND2X1_319 INVX8_23/A INVX1_150/Y gnd NAND2X1_319/Y vdd NAND2X1
XNAND2X1_308 BUFX4_208/Y OAI21X1_699/Y gnd NAND2X1_308/Y vdd NAND2X1
XDFFSR_159 INVX1_52/A CLKBUF1_39/Y DFFSR_167/R vdd DFFSR_159/D gnd vdd DFFSR
XNOR2X1_341 INVX2_43/A INVX4_11/A gnd OAI22X1_43/D vdd NOR2X1
XFILL_21_5_0 gnd vdd FILL
XNOR2X1_330 INVX8_15/A OR2X2_21/B gnd AND2X2_32/A vdd NOR2X1
XFILL_29_6_0 gnd vdd FILL
XFILL_4_6_0 gnd vdd FILL
XFILL_12_5_0 gnd vdd FILL
XNAND3X1_70 wb_adr_i[4] DFFSR_33/Q NOR2X1_3/Y gnd NAND3X1_70/Y vdd NAND3X1
XNAND3X1_92 NAND3X1_92/A NAND3X1_92/B AOI22X1_14/Y gnd DFFSR_87/D vdd NAND3X1
XNAND3X1_81 wb_adr_i[4] INVX1_17/A NOR2X1_3/Y gnd NAND2X1_50/B vdd NAND3X1
XNOR2X1_92 INVX2_74/Y BUFX4_45/Y gnd NOR2X1_92/Y vdd NOR2X1
XNOR2X1_70 INVX2_56/Y BUFX4_44/Y gnd NOR2X1_70/Y vdd NOR2X1
XNOR2X1_81 INVX1_92/Y BUFX4_43/Y gnd NOR2X1_81/Y vdd NOR2X1
XBUFX2_8 BUFX2_8/A gnd ss_pad_o[5] vdd BUFX2
XNAND2X1_138 OR2X2_7/B NAND2X1_138/B gnd AOI21X1_40/B vdd NAND2X1
XNAND2X1_105 XNOR2X1_4/Y NOR2X1_55/B gnd INVX1_85/A vdd NAND2X1
XNAND2X1_149 AND2X2_21/B AND2X2_21/A gnd NAND2X1_149/Y vdd NAND2X1
XNAND2X1_127 NAND2X1_127/A NAND3X1_169/Y gnd DFFSR_244/D vdd NAND2X1
XNAND2X1_3 BUFX4_72/Y wb_dat_i[26] gnd OAI21X1_5/C vdd NAND2X1
XNAND2X1_116 INVX2_82/Y NOR2X1_99/B gnd NAND2X1_116/Y vdd NAND2X1
XNOR2X1_160 INVX2_152/Y NOR2X1_99/B gnd NOR2X1_160/Y vdd NOR2X1
XOAI21X1_611 AOI21X1_212/Y OAI21X1_610/Y NAND2X1_269/Y gnd DFFSR_164/D vdd OAI21X1
XOAI21X1_600 BUFX4_122/Y OAI21X1_599/Y BUFX4_113/Y gnd OAI21X1_601/B vdd OAI21X1
XOAI21X1_644 NOR2X1_294/Y INVX2_144/Y BUFX4_122/Y gnd AOI21X1_241/C vdd OAI21X1
XOAI21X1_633 INVX2_159/Y BUFX4_85/Y NAND2X1_240/Y gnd OAI21X1_634/B vdd OAI21X1
XAOI21X1_8 DFFSR_123/Q AOI21X1_7/B AOI21X1_8/C gnd AOI21X1_8/Y vdd AOI21X1
XNOR2X1_171 INVX2_161/Y BUFX4_42/Y gnd NOR2X1_171/Y vdd NOR2X1
XOAI21X1_655 NOR2X1_297/Y OAI21X1_655/B OAI21X1_655/C gnd DFFSR_146/D vdd OAI21X1
XOAI21X1_666 NOR2X1_306/Y OAI21X1_665/Y OAI21X1_666/C gnd DFFSR_140/D vdd OAI21X1
XOAI21X1_622 BUFX4_62/Y AOI21X1_223/B OAI21X1_622/C gnd OAI21X1_622/Y vdd OAI21X1
XINVX2_8 INVX2_8/A gnd INVX2_8/Y vdd INVX2
XNOR2X1_193 BUFX4_173/Y INVX1_118/A gnd INVX4_7/A vdd NOR2X1
XNOR2X1_182 BUFX4_175/Y AOI21X1_71/C gnd INVX8_14/A vdd NOR2X1
XOAI21X1_688 INVX1_152/Y DFFSR_133/Q BUFX4_113/Y gnd OAI21X1_688/Y vdd OAI21X1
XOAI21X1_677 BUFX4_60/Y NAND2X1_296/Y OAI21X1_677/C gnd OAI21X1_677/Y vdd OAI21X1
XOAI21X1_699 INVX2_87/Y BUFX4_9/Y OAI21X1_699/C gnd OAI21X1_699/Y vdd OAI21X1
XBUFX2_26 BUFX2_26/A gnd ss_pad_o[23] vdd BUFX2
XBUFX2_15 BUFX2_15/A gnd ss_pad_o[12] vdd BUFX2
XINVX1_40 INVX1_40/A gnd INVX1_40/Y vdd INVX1
XINVX1_84 INVX1_84/A gnd INVX1_84/Y vdd INVX1
XINVX1_95 INVX1_95/A gnd INVX1_95/Y vdd INVX1
XINVX1_73 DFFSR_55/Q gnd INVX1_73/Y vdd INVX1
XINVX1_62 INVX1_62/A gnd INVX1_62/Y vdd INVX1
XINVX1_51 INVX1_51/A gnd INVX1_51/Y vdd INVX1
XBUFX2_59 DFFSR_88/Q gnd wb_dat_o[23] vdd BUFX2
XBUFX2_48 BUFX2_48/A gnd wb_dat_o[12] vdd BUFX2
XBUFX2_37 BUFX2_37/A gnd wb_dat_o[1] vdd BUFX2
XNOR2X1_6 NOR2X1_6/A NOR2X1_6/B gnd NOR2X1_6/Y vdd NOR2X1
XFILL_35_4_0 gnd vdd FILL
XAOI21X1_16 INVX1_91/A BUFX4_190/Y AOI21X1_16/C gnd AOI21X1_16/Y vdd AOI21X1
XAOI21X1_38 XNOR2X1_9/A AOI21X1_38/B INVX2_50/Y gnd AOI21X1_38/Y vdd AOI21X1
XAOI21X1_49 AOI21X1_49/A AOI21X1_49/B INVX8_9/Y gnd AOI21X1_49/Y vdd AOI21X1
XAOI21X1_27 AOI21X1_27/A AOI21X1_27/B NOR2X1_46/Y gnd DFFSR_114/D vdd AOI21X1
XFILL_26_4_0 gnd vdd FILL
XOAI22X1_13 BUFX4_78/Y INVX2_14/Y INVX2_36/Y OAI22X1_4/A gnd NOR2X1_9/A vdd OAI22X1
XFILL_1_4_0 gnd vdd FILL
XOAI22X1_35 BUFX4_199/Y INVX2_29/Y INVX8_5/A INVX1_60/Y gnd AOI21X1_15/C vdd OAI22X1
XOAI22X1_24 BUFX4_199/Y INVX2_24/Y OAI22X1_4/C INVX1_49/Y gnd NOR2X1_13/B vdd OAI22X1
XOAI21X1_485 AOI21X1_168/Y OAI21X1_485/B OAI21X1_485/C gnd DFFSR_198/D vdd OAI21X1
XOAI21X1_430 BUFX4_66/Y OR2X2_13/Y AOI21X1_144/Y gnd AOI21X1_146/B vdd OAI21X1
XOAI21X1_474 BUFX4_221/Y OAI21X1_474/B BUFX4_49/Y gnd AOI21X1_166/A vdd OAI21X1
XOAI21X1_441 BUFX4_223/Y OAI21X1_440/Y BUFX4_50/Y gnd OAI21X1_441/Y vdd OAI21X1
XOAI21X1_452 BUFX4_207/Y BUFX4_29/Y INVX2_69/A gnd OAI21X1_452/Y vdd OAI21X1
XOAI21X1_463 BUFX4_168/Y OAI21X1_462/Y BUFX4_38/Y gnd OAI21X1_463/Y vdd OAI21X1
XOAI21X1_496 BUFX4_222/Y OAI21X1_496/B BUFX4_49/Y gnd AOI21X1_173/A vdd OAI21X1
XFILL_9_5_0 gnd vdd FILL
XFILL_17_4_0 gnd vdd FILL
XOAI21X1_90 INVX2_22/Y BUFX4_85/Y OAI21X1_90/C gnd OAI21X1_90/Y vdd OAI21X1
XOAI21X1_271 NOR2X1_176/A NAND2X1_134/Y OAI21X1_271/C gnd NOR2X1_175/B vdd OAI21X1
XOAI21X1_282 INVX1_108/Y AOI21X1_48/B AOI21X1_48/Y gnd NAND2X1_150/B vdd OAI21X1
XOAI21X1_293 INVX2_146/Y BUFX4_172/Y OAI21X1_293/C gnd AOI22X1_37/C vdd OAI21X1
XOAI21X1_260 NOR2X1_164/Y NOR2X1_165/Y BUFX4_188/Y gnd OAI21X1_260/Y vdd OAI21X1
XFILL_36_4 gnd vdd FILL
XFILL_32_2_0 gnd vdd FILL
XFILL_23_2_0 gnd vdd FILL
XDFFSR_82 BUFX2_53/A DFFSR_82/CLK DFFSR_2/R vdd DFFSR_82/D gnd vdd DFFSR
XDFFSR_71 BUFX2_42/A DFFSR_71/CLK DFFSR_2/R vdd DFFSR_71/D gnd vdd DFFSR
XDFFSR_60 INVX2_28/A CLKBUF1_5/A DFFSR_58/R vdd DFFSR_60/D gnd vdd DFFSR
XDFFSR_93 BUFX2_64/A DFFSR_78/CLK DFFSR_95/R vdd DFFSR_93/D gnd vdd DFFSR
XFILL_6_3_0 gnd vdd FILL
XFILL_14_2_0 gnd vdd FILL
XINVX1_132 NOR2X1_19/Y gnd INVX1_132/Y vdd INVX1
XINVX1_110 INVX1_110/A gnd INVX1_110/Y vdd INVX1
XINVX1_143 INVX1_143/A gnd INVX1_143/Y vdd INVX1
XINVX1_154 INVX1_154/A gnd INVX1_154/Y vdd INVX1
XINVX1_121 NOR3X1_3/B gnd INVX1_121/Y vdd INVX1
XAOI21X1_114 BUFX4_151/Y OAI21X1_367/Y BUFX4_47/Y gnd AOI21X1_115/A vdd AOI21X1
XAOI21X1_103 NOR2X1_188/Y BUFX4_65/Y AOI21X1_103/C gnd OAI21X1_320/A vdd AOI21X1
XAOI21X1_169 NOR2X1_252/Y BUFX4_58/Y AOI21X1_169/C gnd AOI21X1_169/Y vdd AOI21X1
XAOI21X1_147 INVX2_104/Y AOI21X1_147/B BUFX4_152/Y gnd OAI21X1_432/C vdd AOI21X1
XAOI21X1_136 NOR2X1_226/Y BUFX4_59/Y AOI21X1_136/C gnd OAI21X1_420/A vdd AOI21X1
XAOI21X1_158 MUX2X1_4/B NAND2X1_250/Y BUFX4_229/Y gnd AOI21X1_158/Y vdd AOI21X1
XAOI21X1_125 BUFX4_148/Y OAI21X1_383/Y BUFX4_49/Y gnd AOI21X1_125/Y vdd AOI21X1
XNAND3X1_129 INVX8_10/Y NAND3X1_129/B OAI21X1_224/Y gnd NAND3X1_129/Y vdd NAND3X1
XNAND3X1_107 INVX1_74/Y AND2X2_4/Y AND2X2_5/Y gnd NOR2X1_44/B vdd NAND3X1
XNAND3X1_118 INVX8_10/A OAI21X1_214/Y NAND3X1_118/C gnd NAND3X1_118/Y vdd NAND3X1
XDFFSR_116 DFFSR_116/Q DFFSR_71/CLK DFFSR_165/R vdd DFFSR_116/D gnd vdd DFFSR
XFILL_30_5_1 gnd vdd FILL
XDFFSR_149 INVX1_29/A CLKBUF1_6/A BUFX4_130/Y vdd DFFSR_149/D gnd vdd DFFSR
XDFFSR_138 INVX2_56/A CLKBUF1_12/Y DFFSR_137/R vdd DFFSR_138/D gnd vdd DFFSR
XDFFSR_105 XNOR2X1_1/B CLKBUF1_38/A vdd BUFX4_87/Y DFFSR_105/D gnd vdd DFFSR
XDFFSR_127 INVX1_97/A CLKBUF1_45/Y DFFSR_130/R vdd DFFSR_127/D gnd vdd DFFSR
XNAND2X1_309 INVX1_156/A BUFX4_62/Y gnd AOI22X1_82/C vdd NAND2X1
XNOR2X1_342 INVX2_48/A INVX4_11/A gnd NOR2X1_342/Y vdd NOR2X1
XNOR2X1_320 INVX1_158/A BUFX4_61/Y gnd NOR2X1_320/Y vdd NOR2X1
XNOR2X1_331 INVX2_130/A BUFX4_37/Y gnd NOR2X1_331/Y vdd NOR2X1
XFILL_21_5_1 gnd vdd FILL
XFILL_20_0_0 gnd vdd FILL
XFILL_29_6_1 gnd vdd FILL
XFILL_28_1_0 gnd vdd FILL
XFILL_4_6_1 gnd vdd FILL
XFILL_3_1_0 gnd vdd FILL
XFILL_11_0_0 gnd vdd FILL
XFILL_12_5_1 gnd vdd FILL
XNOR2X1_60 INVX2_42/A INVX2_49/Y gnd NOR2X1_60/Y vdd NOR2X1
XNAND3X1_71 wb_adr_i[3] INVX2_146/A NOR2X1_4/Y gnd NAND3X1_71/Y vdd NAND3X1
XNAND3X1_60 AND2X2_2/B NAND3X1_60/B BUFX4_107/Y gnd NAND3X1_60/Y vdd NAND3X1
XNAND3X1_93 AOI22X1_16/Y NAND2X1_67/Y AOI22X1_15/Y gnd DFFSR_88/D vdd NAND3X1
XNOR2X1_71 INVX2_57/Y NOR2X1_71/B gnd NOR2X1_71/Y vdd NOR2X1
XFILL_19_1_0 gnd vdd FILL
XNAND3X1_82 wb_adr_i[3] INVX2_72/A NOR2X1_4/Y gnd NAND2X1_52/A vdd NAND3X1
XNOR2X1_82 INVX2_66/Y NOR2X1_99/B gnd NOR2X1_82/Y vdd NOR2X1
XNOR2X1_93 INVX2_75/Y BUFX4_217/Y gnd NOR2X1_93/Y vdd NOR2X1
XBUFX2_9 BUFX2_9/A gnd ss_pad_o[6] vdd BUFX2
XNAND2X1_139 INVX2_43/A INVX2_48/A gnd NOR2X1_176/B vdd NAND2X1
XNAND2X1_106 NAND2X1_106/A INVX1_86/Y gnd INVX1_107/A vdd NAND2X1
XNAND2X1_128 INVX8_13/Y INVX1_89/A gnd AOI22X1_36/A vdd NAND2X1
XNAND2X1_4 MUX2X1_6/S wb_dat_i[27] gnd OAI21X1_7/C vdd NAND2X1
XNAND2X1_117 INVX2_96/Y INVX8_10/A gnd OAI21X1_227/C vdd NAND2X1
XNOR2X1_150 INVX2_144/Y BUFX4_45/Y gnd NOR2X1_150/Y vdd NOR2X1
XNOR2X1_172 INVX2_162/Y NOR2X1_71/B gnd NOR2X1_172/Y vdd NOR2X1
XNOR2X1_183 INVX1_114/A INVX1_113/A gnd INVX2_164/A vdd NOR2X1
XNOR2X1_194 BUFX4_175/Y AOI21X1_69/C gnd INVX8_17/A vdd NOR2X1
XNOR2X1_161 INVX1_101/Y BUFX4_43/Y gnd NOR2X1_161/Y vdd NOR2X1
XINVX2_9 DFFSR_1/Q gnd INVX2_9/Y vdd INVX2
XOAI21X1_601 OAI21X1_601/A OAI21X1_601/B NAND2X1_267/Y gnd DFFSR_166/D vdd OAI21X1
XOAI21X1_645 INVX2_144/Y BUFX4_81/Y NAND2X1_245/Y gnd OAI21X1_645/Y vdd OAI21X1
XOAI21X1_689 NOR2X1_311/Y OAI21X1_688/Y OAI21X1_689/C gnd DFFSR_133/D vdd OAI21X1
XOAI21X1_634 BUFX4_121/Y OAI21X1_634/B BUFX4_114/Y gnd OAI21X1_635/B vdd OAI21X1
XOAI21X1_667 INVX1_149/Y INVX8_22/Y INVX2_56/Y gnd OAI21X1_667/Y vdd OAI21X1
XOAI21X1_678 OAI21X1_677/Y INVX8_21/A OAI21X1_678/C gnd DFFSR_136/D vdd OAI21X1
XAOI21X1_9 INVX2_96/A AOI21X1_7/B AOI21X1_9/C gnd AOI21X1_9/Y vdd AOI21X1
XOAI21X1_656 NOR2X1_1/A INVX8_18/Y NOR2X1_266/Y gnd NOR2X1_316/B vdd OAI21X1
XOAI21X1_623 INVX2_71/Y BUFX4_12/Y NAND2X1_236/Y gnd AOI21X1_224/B vdd OAI21X1
XOAI21X1_612 BUFX4_62/Y NAND2X1_270/Y OAI21X1_612/C gnd AOI21X1_215/B vdd OAI21X1
XBUFX2_38 BUFX2_38/A gnd wb_dat_o[2] vdd BUFX2
XINVX1_85 INVX1_85/A gnd INVX1_85/Y vdd INVX1
XINVX1_30 INVX1_30/A gnd INVX1_30/Y vdd INVX1
XINVX1_41 INVX1_41/A gnd INVX1_41/Y vdd INVX1
XBUFX2_16 BUFX2_16/A gnd ss_pad_o[13] vdd BUFX2
XBUFX2_27 BUFX2_27/A gnd ss_pad_o[24] vdd BUFX2
XINVX1_96 INVX1_96/A gnd INVX1_96/Y vdd INVX1
XINVX1_74 NOR3X1_2/B gnd INVX1_74/Y vdd INVX1
XINVX1_63 INVX1_63/A gnd INVX1_63/Y vdd INVX1
XINVX1_52 INVX1_52/A gnd INVX1_52/Y vdd INVX1
XBUFX2_49 BUFX2_49/A gnd wb_dat_o[13] vdd BUFX2
XNOR2X1_7 NOR2X1_7/A NOR2X1_7/B gnd NOR2X1_7/Y vdd NOR2X1
XFILL_35_4_1 gnd vdd FILL
XAOI21X1_39 AOI21X1_39/A NOR2X1_178/Y AOI21X1_38/Y gnd INVX1_116/A vdd AOI21X1
XAOI21X1_28 INVX1_88/Y AND2X2_10/A NOR2X1_56/Y gnd AND2X2_11/A vdd AOI21X1
XAOI21X1_17 DFFSR_163/Q AOI22X1_7/B OAI22X1_37/Y gnd NAND2X1_59/A vdd AOI21X1
XFILL_26_4_1 gnd vdd FILL
XOAI22X1_14 OAI22X1_4/C INVX1_38/Y INVX1_39/Y INVX8_5/A gnd NOR2X1_9/B vdd OAI22X1
XFILL_1_4_1 gnd vdd FILL
XOAI22X1_25 BUFX4_77/Y INVX2_3/Y INVX1_50/Y BUFX4_226/Y gnd NOR2X1_14/A vdd OAI22X1
XOAI22X1_36 BUFX4_77/Y INVX2_7/Y INVX1_61/Y BUFX4_226/Y gnd AOI21X1_16/C vdd OAI22X1
XOAI21X1_486 BUFX4_211/Y BUFX4_28/Y AOI22X1_3/D gnd OAI21X1_490/C vdd OAI21X1
XOAI21X1_431 INVX2_145/Y BUFX4_82/Y NAND2X1_245/Y gnd OAI21X1_431/Y vdd OAI21X1
XOAI21X1_475 INVX8_21/A BUFX4_31/Y DFFSR_199/Q gnd OAI21X1_475/Y vdd OAI21X1
XOAI21X1_442 BUFX4_207/Y BUFX4_29/Y INVX2_83/A gnd OAI21X1_442/Y vdd OAI21X1
XOAI21X1_453 AND2X2_23/Y INVX2_69/Y BUFX4_168/Y gnd AOI21X1_157/C vdd OAI21X1
XOAI21X1_464 OAI21X1_464/A OAI21X1_463/Y OAI21X1_460/Y gnd DFFSR_204/D vdd OAI21X1
XOAI21X1_497 BUFX4_203/Y BUFX4_30/Y INVX1_58/A gnd OAI21X1_497/Y vdd OAI21X1
XOAI21X1_420 OAI21X1_420/A OAI21X1_420/B OAI21X1_416/Y gnd DFFSR_217/D vdd OAI21X1
XFILL_8_0_0 gnd vdd FILL
XFILL_9_5_1 gnd vdd FILL
XFILL_17_4_1 gnd vdd FILL
XOAI21X1_91 AND2X2_2/Y INVX2_22/Y NAND3X1_48/Y gnd DFFSR_39/D vdd OAI21X1
XOAI21X1_80 INVX1_23/Y BUFX4_80/Y NAND2X1_26/Y gnd NAND3X1_43/A vdd OAI21X1
XOAI21X1_250 NOR2X1_146/Y NOR2X1_147/Y BUFX4_194/Y gnd NAND3X1_152/B vdd OAI21X1
XOAI21X1_272 INVX1_103/A INVX8_13/Y INVX2_48/Y gnd OAI21X1_272/Y vdd OAI21X1
XOAI21X1_283 NAND2X1_104/Y BUFX4_112/Y NAND2X1_134/Y gnd NAND2X1_151/B vdd OAI21X1
XOAI21X1_294 AOI21X1_53/Y INVX1_106/A NAND2X1_149/Y gnd INVX1_118/A vdd OAI21X1
XOAI21X1_261 NOR2X1_166/Y NOR2X1_167/Y BUFX4_184/Y gnd NAND3X1_163/B vdd OAI21X1
XFILL_32_2_1 gnd vdd FILL
XFILL_23_2_1 gnd vdd FILL
XDFFSR_83 DFFSR_83/Q DFFSR_83/CLK DFFSR_88/R vdd DFFSR_83/D gnd vdd DFFSR
XDFFSR_50 OR2X2_2/A DFFSR_5/CLK DFFSR_9/R vdd DFFSR_50/D gnd vdd DFFSR
XDFFSR_72 BUFX2_43/A DFFSR_87/CLK DFFSR_9/R vdd DFFSR_72/D gnd vdd DFFSR
XDFFSR_94 DFFSR_94/Q CLKBUF1_8/Y DFFSR_25/R vdd DFFSR_94/D gnd vdd DFFSR
XDFFSR_61 INVX2_29/A DFFSR_61/CLK DFFSR_95/R vdd DFFSR_61/D gnd vdd DFFSR
XFILL_6_3_1 gnd vdd FILL
XFILL_14_2_1 gnd vdd FILL
XINVX1_100 DFFSR_133/Q gnd INVX1_100/Y vdd INVX1
XINVX1_144 INVX1_144/A gnd INVX1_144/Y vdd INVX1
XINVX1_133 INVX1_133/A gnd INVX1_133/Y vdd INVX1
XINVX1_111 INVX1_111/A gnd INVX1_111/Y vdd INVX1
XINVX1_122 INVX1_122/A gnd INVX1_122/Y vdd INVX1
XINVX1_155 INVX1_155/A gnd INVX1_155/Y vdd INVX1
XFILL_27_1 gnd vdd FILL
XAOI21X1_115 AOI21X1_115/A OAI21X1_366/Y NOR2X1_213/Y gnd DFFSR_232/D vdd AOI21X1
XAOI21X1_148 BUFX4_151/Y OAI21X1_433/Y BUFX4_48/Y gnd AOI21X1_149/A vdd AOI21X1
XAOI21X1_137 INVX2_93/Y AOI21X1_137/B BUFX4_150/Y gnd OAI21X1_421/C vdd AOI21X1
XAOI21X1_104 AND2X2_22/Y BUFX4_65/Y OAI21X1_322/Y gnd OAI21X1_325/A vdd AOI21X1
XAOI21X1_126 AOI21X1_125/Y AOI21X1_126/B NOR2X1_218/Y gnd DFFSR_226/D vdd AOI21X1
XAOI21X1_159 AOI21X1_159/A AOI21X1_159/B NOR2X1_240/Y gnd DFFSR_205/D vdd AOI21X1
XNAND3X1_108 BUFX4_245/Y NAND3X1_108/B OR2X2_9/Y gnd OAI21X1_203/C vdd NAND3X1
XNAND3X1_119 INVX4_4/Y NAND3X1_117/Y NAND3X1_118/Y gnd NAND3X1_119/Y vdd NAND3X1
XDFFSR_117 INVX1_99/A CLKBUF1_27/Y DFFSR_165/R vdd DFFSR_117/D gnd vdd DFFSR
XDFFSR_139 DFFSR_139/Q CLKBUF1_5/Y DFFSR_151/R vdd DFFSR_139/D gnd vdd DFFSR
XDFFSR_128 INVX2_87/A DFFSR_8/CLK DFFSR_151/R vdd DFFSR_128/D gnd vdd DFFSR
XDFFSR_106 DFFSR_106/Q DFFSR_61/CLK vdd BUFX4_87/Y DFFSR_106/D gnd vdd DFFSR
XNOR2X1_343 INVX4_11/Y INVX1_90/A gnd OAI22X1_45/C vdd NOR2X1
XNOR2X1_310 BUFX4_28/Y NOR2X1_310/B gnd NOR2X1_310/Y vdd NOR2X1
XNOR2X1_321 NOR2X1_321/A BUFX4_64/Y gnd NOR2X1_321/Y vdd NOR2X1
XNOR2X1_332 INVX8_22/Y NOR2X1_337/B gnd INVX1_162/A vdd NOR2X1
XFILL_20_0_1 gnd vdd FILL
XFILL_28_1_1 gnd vdd FILL
XFILL_3_1_1 gnd vdd FILL
XFILL_11_0_1 gnd vdd FILL
XNAND3X1_50 wb_adr_i[4] wb_adr_i[2] INVX2_17/Y gnd BUFX4_200/A vdd NAND3X1
XNOR2X1_61 INVX2_49/A INVX2_42/Y gnd NOR2X1_62/B vdd NOR2X1
XNOR2X1_50 NOR2X1_50/A INVX1_79/Y gnd OR2X2_3/B vdd NOR2X1
XNAND3X1_72 wb_adr_i[4] INVX2_46/A NOR2X1_3/Y gnd NAND3X1_72/Y vdd NAND3X1
XNAND3X1_61 BUFX4_15/Y NAND3X1_61/B BUFX4_107/Y gnd NAND3X1_61/Y vdd NAND3X1
XNOR2X1_94 INVX2_76/Y BUFX4_44/Y gnd NOR2X1_94/Y vdd NOR2X1
XNOR2X1_72 INVX2_58/Y BUFX4_44/Y gnd NOR2X1_72/Y vdd NOR2X1
XFILL_19_1_1 gnd vdd FILL
XNAND3X1_83 wb_adr_i[4] DFFSR_43/Q NOR2X1_3/Y gnd NAND2X1_52/B vdd NAND3X1
XNAND3X1_94 NAND3X1_94/A NAND3X1_94/B NAND3X1_94/C gnd DFFSR_89/D vdd NAND3X1
XNOR2X1_83 INVX2_67/Y NOR2X1_87/B gnd NOR2X1_83/Y vdd NOR2X1
XNAND2X1_107 AOI21X1_46/A OR2X2_7/A gnd NAND2X1_107/Y vdd NAND2X1
XNAND2X1_129 NAND2X1_129/A NAND2X1_129/B gnd NOR2X1_180/B vdd NAND2X1
XNAND2X1_5 MUX2X1_8/S wb_dat_i[28] gnd OAI21X1_9/C vdd NAND2X1
XNAND2X1_118 INVX2_97/Y BUFX4_238/Y gnd OAI21X1_228/C vdd NAND2X1
XNOR2X1_184 DFFSR_33/Q INVX8_9/Y gnd XOR2X1_4/B vdd NOR2X1
XNOR2X1_151 INVX2_145/Y BUFX4_217/Y gnd NOR2X1_151/Y vdd NOR2X1
XNOR2X1_173 INVX2_163/Y BUFX4_42/Y gnd NOR2X1_173/Y vdd NOR2X1
XNOR2X1_195 BUFX4_155/Y AOI21X1_71/C gnd INVX4_9/A vdd NOR2X1
XNOR2X1_162 INVX2_153/Y NOR2X1_76/B gnd NOR2X1_162/Y vdd NOR2X1
XNOR2X1_140 INVX2_126/Y BUFX4_43/Y gnd NOR2X1_140/Y vdd NOR2X1
XOAI21X1_646 BUFX4_122/Y OAI21X1_645/Y BUFX4_113/Y gnd OAI21X1_646/Y vdd OAI21X1
XOAI21X1_602 BUFX4_101/Y INVX8_11/Y INVX1_137/A gnd NOR2X1_310/B vdd OAI21X1
XOAI21X1_635 OAI21X1_635/A OAI21X1_635/B NAND2X1_277/Y gnd DFFSR_153/D vdd OAI21X1
XOAI21X1_668 BUFX4_58/Y NAND2X1_290/Y OAI21X1_667/Y gnd OAI21X1_668/Y vdd OAI21X1
XOAI21X1_679 INVX2_119/Y BUFX4_164/Y NAND2X1_222/Y gnd NAND2X1_297/B vdd OAI21X1
XOAI21X1_657 NOR2X1_1/A INVX8_18/Y AND2X2_30/A gnd OR2X2_18/A vdd OAI21X1
XOAI21X1_613 INVX2_61/Y BUFX4_8/Y NAND2X1_231/Y gnd AOI21X1_214/B vdd OAI21X1
XOAI21X1_624 NOR2X1_287/Y MUX2X1_1/A BUFX4_120/Y gnd AOI21X1_226/C vdd OAI21X1
XINVX1_31 INVX1_31/A gnd INVX1_31/Y vdd INVX1
XINVX1_42 INVX1_42/A gnd INVX1_42/Y vdd INVX1
XINVX1_20 DFFSR_41/Q gnd INVX1_20/Y vdd INVX1
XINVX1_86 INVX1_86/A gnd INVX1_86/Y vdd INVX1
XBUFX2_39 DFFSR_68/Q gnd wb_dat_o[3] vdd BUFX2
XINVX1_64 DFFSR_63/Q gnd INVX1_64/Y vdd INVX1
XBUFX2_17 BUFX2_17/A gnd ss_pad_o[14] vdd BUFX2
XBUFX2_28 BUFX2_28/A gnd ss_pad_o[25] vdd BUFX2
XINVX1_75 INVX1_75/A gnd INVX1_75/Y vdd INVX1
XINVX1_97 INVX1_97/A gnd INVX1_97/Y vdd INVX1
XINVX1_53 INVX1_53/A gnd INVX1_53/Y vdd INVX1
XNOR2X1_8 NOR2X1_8/A NOR2X1_8/B gnd NOR2X1_8/Y vdd NOR2X1
XAOI21X1_29 NOR2X1_60/Y XOR2X1_2/B NOR2X1_65/Y gnd AOI21X1_29/Y vdd AOI21X1
XAOI21X1_18 INVX1_98/A BUFX4_190/Y AOI21X1_18/C gnd NAND2X1_59/B vdd AOI21X1
XOAI22X1_15 OAI22X1_9/A INVX1_40/Y INVX8_2/A INVX2_21/Y gnd AOI21X1_6/C vdd OAI22X1
XOAI21X1_432 BUFX4_66/Y AOI21X1_147/B OAI21X1_432/C gnd AOI21X1_149/B vdd OAI21X1
XOAI21X1_421 BUFX4_60/Y AOI21X1_137/B OAI21X1_421/C gnd OAI21X1_421/Y vdd OAI21X1
XOAI22X1_37 BUFX4_199/Y INVX2_30/Y INVX1_62/Y BUFX4_226/Y gnd OAI22X1_37/Y vdd OAI22X1
XOAI22X1_26 BUFX4_199/Y INVX2_25/Y OAI22X1_4/C INVX1_51/Y gnd NOR2X1_14/B vdd OAI22X1
XOAI21X1_410 OAI21X1_410/A OAI21X1_410/B OAI21X1_410/C gnd DFFSR_220/D vdd OAI21X1
XOAI21X1_487 NOR2X1_252/Y INVX2_149/Y BUFX4_171/Y gnd AOI21X1_169/C vdd OAI21X1
XOAI21X1_465 BUFX4_66/Y OAI21X1_465/B AOI21X1_161/Y gnd OAI21X1_465/Y vdd OAI21X1
XOAI21X1_476 BUFX4_98/Y INVX4_6/Y INVX1_128/Y gnd NOR2X1_262/B vdd OAI21X1
XOAI21X1_454 INVX2_69/Y MUX2X1_8/S OAI21X1_572/C gnd OAI21X1_455/B vdd OAI21X1
XOAI21X1_498 NOR2X1_256/Y INVX2_155/Y BUFX4_167/Y gnd AOI21X1_174/C vdd OAI21X1
XOAI21X1_443 BUFX4_99/Y INVX4_6/Y INVX1_124/A gnd NOR2X1_257/B vdd OAI21X1
XFILL_8_0_1 gnd vdd FILL
XOAI21X1_81 AND2X2_2/Y INVX1_23/Y OAI21X1_81/C gnd DFFSR_34/D vdd OAI21X1
XOAI21X1_70 AND2X2_2/Y INVX2_18/Y NAND3X1_38/Y gnd DFFSR_44/D vdd OAI21X1
XOAI21X1_92 INVX1_25/Y BUFX4_86/Y OAI21X1_92/C gnd OAI21X1_92/Y vdd OAI21X1
XOAI21X1_273 AOI21X1_34/Y OAI21X1_273/B AOI21X1_35/Y gnd NAND2X1_144/B vdd OAI21X1
XOAI21X1_262 NOR2X1_168/Y NOR2X1_169/Y BUFX4_194/Y gnd OAI21X1_262/Y vdd OAI21X1
XOAI21X1_251 NOR2X1_148/Y NOR2X1_149/Y BUFX4_185/Y gnd NAND3X1_152/C vdd OAI21X1
XOAI21X1_240 NOR2X1_127/Y NOR2X1_128/Y BUFX4_194/Y gnd OAI21X1_240/Y vdd OAI21X1
XFILL_10_6_0 gnd vdd FILL
XOAI21X1_284 XNOR2X1_11/Y INVX8_9/Y OAI21X1_284/C gnd INVX1_114/A vdd OAI21X1
XOAI21X1_295 INVX2_149/Y BUFX4_172/Y OAI21X1_295/C gnd AOI22X1_38/C vdd OAI21X1
XNAND2X1_290 INVX8_22/A INVX1_149/A gnd NAND2X1_290/Y vdd NAND2X1
XDFFSR_40 DFFSR_40/Q DFFSR_85/CLK DFFSR_1/R vdd DFFSR_40/D gnd vdd DFFSR
XDFFSR_51 DFFSR_51/Q DFFSR_6/CLK DFFSR_7/R vdd DFFSR_51/D gnd vdd DFFSR
XDFFSR_84 BUFX2_55/A DFFSR_9/CLK DFFSR_9/R vdd DFFSR_84/D gnd vdd DFFSR
XDFFSR_73 BUFX2_44/A CLKBUF1_23/Y DFFSR_53/R vdd DFFSR_73/D gnd vdd DFFSR
XDFFSR_95 BUFX2_66/A CLKBUF1_2/Y DFFSR_95/R vdd DFFSR_95/D gnd vdd DFFSR
XDFFSR_62 INVX2_30/A DFFSR_47/CLK DFFSR_58/R vdd DFFSR_62/D gnd vdd DFFSR
XCLKBUF1_60 wb_clk_i gnd CLKBUF1_8/A vdd CLKBUF1
XINVX1_101 MUX2X1_5/B gnd INVX1_101/Y vdd INVX1
XINVX1_112 INVX1_112/A gnd INVX1_112/Y vdd INVX1
XINVX1_134 INVX1_134/A gnd INVX1_134/Y vdd INVX1
XINVX1_123 INVX1_123/A gnd INVX1_123/Y vdd INVX1
XINVX1_145 INVX1_145/A gnd INVX1_145/Y vdd INVX1
XINVX1_156 INVX1_156/A gnd INVX1_156/Y vdd INVX1
XFILL_33_5_0 gnd vdd FILL
XFILL_27_2 gnd vdd FILL
XAOI21X1_149 AOI21X1_149/A AOI21X1_149/B NOR2X1_231/Y gnd DFFSR_212/D vdd AOI21X1
XAOI21X1_138 BUFX4_150/Y OAI21X1_422/Y BUFX4_48/Y gnd AOI21X1_139/A vdd AOI21X1
XAOI21X1_116 INVX2_120/Y NAND2X1_221/Y INVX8_15/A gnd OAI21X1_368/C vdd AOI21X1
XAOI21X1_105 NOR2X1_204/Y BUFX4_65/Y AOI21X1_105/C gnd OAI21X1_330/A vdd AOI21X1
XAOI21X1_127 NOR2X1_219/Y BUFX4_67/Y AOI21X1_127/C gnd OAI21X1_388/A vdd AOI21X1
XFILL_24_5_0 gnd vdd FILL
XNAND3X1_109 BUFX4_194/Y NAND2X1_111/Y NAND3X1_109/C gnd NAND3X1_110/B vdd NAND3X1
XFILL_7_6_0 gnd vdd FILL
XFILL_15_5_0 gnd vdd FILL
XDFFSR_107 DFFSR_107/Q DFFSR_47/CLK vdd BUFX4_90/Y DFFSR_107/D gnd vdd DFFSR
XDFFSR_118 INVX2_74/A CLKBUF1_23/Y DFFSR_137/R vdd DFFSR_118/D gnd vdd DFFSR
XDFFSR_129 DFFSR_129/Q DFFSR_99/CLK DFFSR_130/R vdd DFFSR_129/D gnd vdd DFFSR
XBUFX4_240 INVX8_16/Y gnd BUFX4_240/Y vdd BUFX4
XNOR2X1_344 XOR2X1_3/B INVX4_5/A gnd AND2X2_33/A vdd NOR2X1
XNOR2X1_311 INVX1_152/A BUFX4_61/Y gnd NOR2X1_311/Y vdd NOR2X1
XNOR2X1_322 INVX1_159/A BUFX4_58/Y gnd NOR2X1_322/Y vdd NOR2X1
XNOR2X1_300 INVX8_22/Y NOR2X1_300/B gnd INVX1_144/A vdd NOR2X1
XNOR2X1_333 DFFSR_163/Q BUFX4_118/Y gnd NOR2X1_333/Y vdd NOR2X1
XNAND3X1_73 wb_adr_i[3] INVX2_73/A NOR2X1_4/Y gnd NAND3X1_73/Y vdd NAND3X1
XNAND3X1_62 AND2X2_2/B NAND3X1_62/B BUFX4_106/Y gnd NAND3X1_62/Y vdd NAND3X1
XNAND3X1_40 OAI21X1_73/Y BUFX4_18/Y INVX8_2/Y gnd OAI21X1_74/C vdd NAND3X1
XNAND3X1_51 BUFX4_20/Y NAND3X1_51/B AND2X2_3/A gnd OAI21X1_95/C vdd NAND3X1
XNAND3X1_84 wb_adr_i[3] INVX2_86/A NOR2X1_4/Y gnd NAND3X1_84/Y vdd NAND3X1
XNOR2X1_62 NOR2X1_60/Y NOR2X1_62/B gnd INVX1_87/A vdd NOR2X1
XNOR2X1_73 INVX2_59/Y NOR2X1_97/B gnd NOR2X1_73/Y vdd NOR2X1
XNOR2X1_95 INVX2_77/Y NOR2X1_97/B gnd NOR2X1_95/Y vdd NOR2X1
XNOR2X1_51 NOR2X1_51/A OR2X2_3/B gnd NOR2X1_51/Y vdd NOR2X1
XNAND3X1_95 NAND3X1_95/A NAND3X1_95/B NAND3X1_95/C gnd DFFSR_90/D vdd NAND3X1
XNOR2X1_40 NOR3X1_2/A NOR3X1_2/C gnd NOR2X1_40/Y vdd NOR2X1
XNOR2X1_84 INVX2_68/Y BUFX4_40/Y gnd NOR2X1_84/Y vdd NOR2X1
XFILL_30_3_0 gnd vdd FILL
XNAND2X1_108 NAND2X1_108/A OR2X2_7/Y gnd INVX1_90/A vdd NAND2X1
XNAND2X1_119 INVX2_98/Y BUFX4_238/Y gnd OAI21X1_230/C vdd NAND2X1
XNAND2X1_6 BUFX4_71/Y wb_dat_i[29] gnd NAND2X1_6/Y vdd NAND2X1
XNOR2X1_163 INVX2_154/Y BUFX4_41/Y gnd NOR2X1_163/Y vdd NOR2X1
XOAI21X1_603 NOR2X1_281/Y INVX2_147/Y BUFX4_121/Y gnd AOI21X1_211/C vdd OAI21X1
XNOR2X1_152 INVX1_99/Y BUFX4_45/Y gnd NOR2X1_152/Y vdd NOR2X1
XFILL_21_3_0 gnd vdd FILL
XNOR2X1_130 INVX2_117/Y BUFX4_46/Y gnd NOR2X1_130/Y vdd NOR2X1
XNOR2X1_185 AOI21X1_50/Y AOI21X1_49/Y gnd INVX1_110/A vdd NOR2X1
XNOR2X1_141 INVX2_127/Y NOR2X1_87/B gnd NOR2X1_141/Y vdd NOR2X1
XNOR2X1_174 BUFX4_99/Y INVX8_11/Y gnd BUFX4_230/A vdd NOR2X1
XOAI21X1_614 BUFX4_64/Y AOI21X1_216/B OAI21X1_614/C gnd AOI21X1_218/B vdd OAI21X1
XNOR2X1_196 BUFX4_155/Y INVX1_117/A gnd INVX8_23/A vdd NOR2X1
XOAI21X1_647 AOI21X1_241/Y OAI21X1_646/Y OAI21X1_647/C gnd DFFSR_149/D vdd OAI21X1
XOAI21X1_669 INVX2_56/Y BUFX4_161/Y OAI21X1_587/C gnd NAND2X1_291/B vdd OAI21X1
XOAI21X1_636 BUFX4_60/Y AOI21X1_234/B OAI21X1_636/C gnd OAI21X1_636/Y vdd OAI21X1
XOAI21X1_658 BUFX4_96/Y INVX8_18/Y AND2X2_29/A gnd NOR2X1_300/B vdd OAI21X1
XOAI21X1_625 MUX2X1_1/A BUFX4_5/Y OAI21X1_515/C gnd OAI21X1_626/B vdd OAI21X1
XINVX1_21 INVX4_11/A gnd INVX1_21/Y vdd INVX1
XINVX1_10 INVX1_10/A gnd INVX1_10/Y vdd INVX1
XINVX1_32 INVX1_32/A gnd INVX1_32/Y vdd INVX1
XINVX1_43 INVX1_43/A gnd INVX1_43/Y vdd INVX1
XINVX1_76 OR2X2_4/A gnd INVX1_76/Y vdd INVX1
XINVX1_65 XOR2X1_1/B gnd INVX1_65/Y vdd INVX1
XINVX1_54 INVX1_54/A gnd INVX1_54/Y vdd INVX1
XINVX1_87 INVX1_87/A gnd INVX1_87/Y vdd INVX1
XFILL_29_4_0 gnd vdd FILL
XBUFX2_29 BUFX2_29/A gnd ss_pad_o[26] vdd BUFX2
XFILL_4_4_0 gnd vdd FILL
XINVX1_98 INVX1_98/A gnd INVX1_98/Y vdd INVX1
XBUFX2_18 BUFX2_18/A gnd ss_pad_o[15] vdd BUFX2
XFILL_12_3_0 gnd vdd FILL
XNOR2X1_9 NOR2X1_9/A NOR2X1_9/B gnd NOR2X1_9/Y vdd NOR2X1
XAOI21X1_19 DFFSR_41/Q OR2X2_1/A BUFX2_2/A gnd OAI22X1_40/D vdd AOI21X1
XOAI21X1_466 INVX2_55/Y BUFX4_161/Y OAI21X1_587/C gnd OAI21X1_466/Y vdd OAI21X1
XOAI21X1_433 INVX2_104/Y BUFX4_84/Y OAI21X1_732/C gnd OAI21X1_433/Y vdd OAI21X1
XOAI22X1_16 INVX8_1/A INVX2_15/Y INVX2_37/Y OAI22X1_7/D gnd NOR2X1_10/A vdd OAI22X1
XOAI21X1_422 INVX2_93/Y BUFX4_84/Y NAND2X1_242/Y gnd OAI21X1_422/Y vdd OAI21X1
XOAI21X1_411 BUFX4_220/Y INVX8_19/A INVX1_43/A gnd OAI21X1_411/Y vdd OAI21X1
XOAI22X1_27 BUFX4_76/Y INVX2_4/Y INVX2_26/Y INVX8_4/A gnd NOR2X1_15/A vdd OAI22X1
XOAI21X1_444 NOR2X1_236/Y INVX2_83/Y BUFX4_168/Y gnd AOI21X1_154/C vdd OAI21X1
XOAI21X1_455 BUFX4_168/Y OAI21X1_455/B BUFX4_35/Y gnd OAI21X1_456/B vdd OAI21X1
XOAI21X1_400 OAI21X1_400/A OAI21X1_399/Y OAI21X1_400/C gnd DFFSR_222/D vdd OAI21X1
XOAI22X1_38 BUFX4_77/Y INVX2_8/Y INVX8_5/A INVX1_63/Y gnd AOI21X1_18/C vdd OAI22X1
XOAI21X1_488 INVX2_149/Y NAND2X1_9/B NAND2X1_226/Y gnd OAI21X1_489/B vdd OAI21X1
XOAI21X1_477 NOR2X1_248/Y INVX2_118/Y BUFX4_166/Y gnd AOI21X1_167/C vdd OAI21X1
XOAI21X1_499 INVX2_155/Y BUFX4_10/Y NAND2X1_232/Y gnd OAI21X1_500/B vdd OAI21X1
XFILL_35_2_0 gnd vdd FILL
XOAI21X1_60 BUFX4_181/Y INVX2_14/Y OAI21X1_60/C gnd DFFSR_6/D vdd OAI21X1
XOAI21X1_82 INVX1_24/Y BUFX4_81/Y NAND2X1_27/Y gnd NAND3X1_44/A vdd OAI21X1
XOAI21X1_93 AND2X2_2/Y INVX1_25/Y OAI21X1_93/C gnd DFFSR_40/D vdd OAI21X1
XOAI21X1_71 INVX1_19/Y BUFX4_8/Y OAI21X1_71/C gnd OAI21X1_71/Y vdd OAI21X1
XFILL_26_2_0 gnd vdd FILL
XFILL_1_2_0 gnd vdd FILL
XOAI21X1_274 NOR2X1_177/Y AOI21X1_36/Y INVX2_49/A gnd AND2X2_20/A vdd OAI21X1
XOAI21X1_285 AOI21X1_44/Y AOI21X1_33/Y NOR2X1_181/Y gnd AOI21X1_49/B vdd OAI21X1
XOAI21X1_296 INVX2_157/Y BUFX4_178/Y OAI21X1_296/C gnd AOI22X1_42/C vdd OAI21X1
XOAI21X1_263 NOR2X1_170/Y NOR2X1_171/Y BUFX4_185/Y gnd OAI21X1_263/Y vdd OAI21X1
XOAI21X1_241 NOR2X1_129/Y NOR2X1_130/Y BUFX4_185/Y gnd NAND3X1_144/C vdd OAI21X1
XFILL_10_6_1 gnd vdd FILL
XOAI21X1_230 DFFSR_204/Q BUFX4_238/Y OAI21X1_230/C gnd AND2X2_15/A vdd OAI21X1
XOAI21X1_252 AOI21X1_30/Y AOI21X1_31/Y INVX4_4/Y gnd OAI21X1_252/Y vdd OAI21X1
XFILL_9_3_0 gnd vdd FILL
XAND2X2_30 AND2X2_30/A INVX4_10/A gnd AND2X2_30/Y vdd AND2X2
XNAND2X1_280 INVX1_31/A BUFX4_211/Y gnd NAND2X1_280/Y vdd NAND2X1
XNAND2X1_291 BUFX4_206/Y NAND2X1_291/B gnd OAI21X1_670/C vdd NAND2X1
XFILL_17_2_0 gnd vdd FILL
XDFFSR_30 INVX1_6/A CLKBUF1_34/A DFFSR_25/R vdd DFFSR_30/D gnd vdd DFFSR
XDFFSR_85 DFFSR_85/Q DFFSR_85/CLK DFFSR_88/R vdd DFFSR_85/D gnd vdd DFFSR
XDFFSR_41 DFFSR_41/Q DFFSR_71/CLK DFFSR_2/R vdd DFFSR_41/D gnd vdd DFFSR
XDFFSR_63 DFFSR_63/Q DFFSR_3/CLK DFFSR_7/R vdd DFFSR_63/D gnd vdd DFFSR
XDFFSR_52 INVX2_36/A DFFSR_7/CLK DFFSR_9/R vdd DFFSR_52/D gnd vdd DFFSR
XDFFSR_74 DFFSR_74/Q CLKBUF1_55/Y DFFSR_53/R vdd DFFSR_74/D gnd vdd DFFSR
XDFFSR_96 BUFX2_67/A CLKBUF1_52/Y DFFSR_95/R vdd DFFSR_96/D gnd vdd DFFSR
XCLKBUF1_61 wb_clk_i gnd CLKBUF1_3/A vdd CLKBUF1
XCLKBUF1_50 CLKBUF1_5/A gnd CLKBUF1_50/Y vdd CLKBUF1
XINVX1_102 DFFSR_121/Q gnd INVX1_102/Y vdd INVX1
XINVX1_113 INVX1_113/A gnd INVX1_113/Y vdd INVX1
XINVX1_135 DFFSR_204/Q gnd INVX1_135/Y vdd INVX1
XINVX1_157 INVX1_157/A gnd INVX1_157/Y vdd INVX1
XINVX1_146 INVX1_146/A gnd INVX1_146/Y vdd INVX1
XINVX1_124 INVX1_124/A gnd INVX1_124/Y vdd INVX1
XFILL_33_5_1 gnd vdd FILL
XFILL_27_3 gnd vdd FILL
XFILL_32_0_0 gnd vdd FILL
XAOI21X1_139 AOI21X1_139/A OAI21X1_421/Y NOR2X1_227/Y gnd DFFSR_216/D vdd AOI21X1
XAOI21X1_117 BUFX4_150/Y AOI21X1_117/B BUFX4_48/Y gnd AOI21X1_118/A vdd AOI21X1
XAOI21X1_106 NOR2X1_206/Y BUFX4_67/Y AOI21X1_106/C gnd OAI21X1_335/A vdd AOI21X1
XAOI21X1_128 NOR2X1_220/Y BUFX4_67/Y OAI21X1_390/Y gnd OAI21X1_393/A vdd AOI21X1
XFILL_24_5_1 gnd vdd FILL
XFILL_23_0_0 gnd vdd FILL
XINVX4_10 INVX4_10/A gnd OR2X2_17/B vdd INVX4
XFILL_6_1_0 gnd vdd FILL
XFILL_7_6_1 gnd vdd FILL
XFILL_15_5_1 gnd vdd FILL
XDFFSR_119 AOI21X1_4/A CLKBUF1_5/A DFFSR_151/R vdd DFFSR_119/D gnd vdd DFFSR
XDFFSR_108 NOR3X1_2/B DFFSR_78/CLK vdd BUFX4_87/Y DFFSR_108/D gnd vdd DFFSR
XFILL_14_0_0 gnd vdd FILL
XBUFX4_241 INVX8_16/Y gnd BUFX4_241/Y vdd BUFX4
XBUFX4_230 BUFX4_230/A gnd BUFX4_230/Y vdd BUFX4
XNOR2X1_301 INVX8_22/Y NOR2X1_301/B gnd INVX1_145/A vdd NOR2X1
XNOR2X1_345 INVX4_11/Y INVX1_79/Y gnd AOI22X1_85/C vdd NOR2X1
XNOR2X1_323 INVX1_160/A BUFX4_61/Y gnd NOR2X1_323/Y vdd NOR2X1
XFILL_32_1 gnd vdd FILL
XNOR2X1_312 BUFX4_28/Y NOR2X1_282/B gnd NOR2X1_312/Y vdd NOR2X1
XNOR2X1_334 INVX2_129/A BUFX4_115/Y gnd NOR2X1_334/Y vdd NOR2X1
XNAND3X1_74 wb_adr_i[4] INVX4_2/A NOR2X1_3/Y gnd NAND2X1_40/B vdd NAND3X1
XNAND3X1_63 BUFX4_15/Y NAND3X1_63/B BUFX4_107/Y gnd NAND3X1_63/Y vdd NAND3X1
XNAND3X1_41 OAI21X1_75/Y BUFX4_15/Y INVX8_2/Y gnd NAND3X1_41/Y vdd NAND3X1
XNAND3X1_30 AND2X2_2/B NAND3X1_30/B BUFX4_27/Y gnd OAI21X1_56/C vdd NAND3X1
XNAND3X1_85 wb_adr_i[4] INVX1_19/A NOR2X1_3/Y gnd NAND2X1_55/B vdd NAND3X1
XNAND3X1_96 NAND3X1_96/A NAND3X1_96/B NAND3X1_96/C gnd DFFSR_91/D vdd NAND3X1
XNOR2X1_30 DFFSR_103/Q INVX1_70/A gnd AND2X2_5/A vdd NOR2X1
XNAND3X1_52 AND2X2_1/B NAND3X1_52/B BUFX4_108/Y gnd OAI21X1_97/C vdd NAND3X1
XNOR2X1_63 INVX1_87/Y AND2X2_11/A gnd NOR2X1_63/Y vdd NOR2X1
XNOR2X1_52 DFFSR_33/Q INVX2_44/Y gnd INVX1_81/A vdd NOR2X1
XNOR2X1_96 INVX2_78/Y BUFX4_44/Y gnd NOR2X1_96/Y vdd NOR2X1
XNOR2X1_74 INVX2_60/Y BUFX4_44/Y gnd NOR2X1_74/Y vdd NOR2X1
XNOR2X1_41 INVX1_72/A NOR3X1_2/C gnd NOR2X1_41/Y vdd NOR2X1
XNOR2X1_85 INVX2_69/Y NOR2X1_87/B gnd NOR2X1_85/Y vdd NOR2X1
XFILL_30_3_1 gnd vdd FILL
XNAND2X1_109 INVX8_9/Y INVX1_90/A gnd OAI21X1_199/C vdd NAND2X1
XNAND2X1_7 BUFX4_73/Y wb_dat_i[30] gnd NAND2X1_7/Y vdd NAND2X1
XNOR2X1_131 INVX2_118/Y BUFX4_215/Y gnd NOR2X1_131/Y vdd NOR2X1
XNOR2X1_142 INVX2_128/Y BUFX4_215/Y gnd NOR2X1_142/Y vdd NOR2X1
XNOR2X1_120 INVX2_109/Y BUFX4_43/Y gnd NOR2X1_120/Y vdd NOR2X1
XNOR2X1_175 INVX4_2/Y NOR2X1_175/B gnd AOI21X1_43/B vdd NOR2X1
XOAI21X1_648 NOR2X1_295/Y INVX2_105/Y BUFX4_122/Y gnd AOI21X1_242/C vdd OAI21X1
XOAI21X1_604 INVX2_147/Y NAND2X1_9/B NAND2X1_226/Y gnd OAI21X1_604/Y vdd OAI21X1
XNOR2X1_153 INVX2_146/Y BUFX4_217/Y gnd NOR2X1_153/Y vdd NOR2X1
XFILL_21_3_1 gnd vdd FILL
XOAI21X1_637 INVX2_92/Y BUFX4_86/Y NAND2X1_242/Y gnd OAI21X1_637/Y vdd OAI21X1
XNOR2X1_186 INVX1_109/Y INVX1_110/Y gnd INVX1_111/A vdd NOR2X1
XOAI21X1_615 INVX2_154/Y BUFX4_9/Y NAND2X1_232/Y gnd AOI21X1_217/B vdd OAI21X1
XOAI21X1_626 BUFX4_120/Y OAI21X1_626/B BUFX4_118/Y gnd OAI21X1_626/Y vdd OAI21X1
XNOR2X1_164 INVX2_155/Y NOR2X1_76/B gnd NOR2X1_164/Y vdd NOR2X1
XNOR2X1_197 BUFX4_173/Y INVX1_117/A gnd INVX4_8/A vdd NOR2X1
XOAI21X1_659 BUFX4_96/Y INVX8_18/Y INVX1_139/Y gnd NOR2X1_301/B vdd OAI21X1
XINVX1_88 INVX1_88/A gnd INVX1_88/Y vdd INVX1
XFILL_29_4_1 gnd vdd FILL
XINVX1_11 INVX1_11/A gnd INVX1_11/Y vdd INVX1
XINVX1_99 INVX1_99/A gnd INVX1_99/Y vdd INVX1
XINVX1_22 DFFSR_33/Q gnd INVX1_22/Y vdd INVX1
XINVX1_33 INVX1_33/A gnd INVX1_33/Y vdd INVX1
XINVX1_44 INVX1_44/A gnd INVX1_44/Y vdd INVX1
XINVX1_55 INVX1_55/A gnd INVX1_55/Y vdd INVX1
XFILL_4_4_1 gnd vdd FILL
XINVX1_77 INVX1_77/A gnd INVX1_77/Y vdd INVX1
XINVX1_66 INVX2_27/A gnd INVX1_66/Y vdd INVX1
XBUFX2_19 BUFX2_19/A gnd ss_pad_o[16] vdd BUFX2
XFILL_12_3_1 gnd vdd FILL
XOAI22X1_39 BUFX2_35/A INVX1_64/Y NAND2X1_33/Y OAI22X1_39/D gnd DFFSR_63/D vdd OAI22X1
XOAI22X1_17 OAI22X1_4/C INVX1_41/Y INVX1_42/Y INVX8_5/A gnd NOR2X1_10/B vdd OAI22X1
XOAI22X1_28 OAI22X1_4/C INVX1_52/Y INVX1_53/Y INVX8_5/A gnd NOR2X1_15/B vdd OAI22X1
XOAI21X1_489 BUFX4_171/Y OAI21X1_489/B BUFX4_36/Y gnd OAI21X1_490/B vdd OAI21X1
XOAI21X1_467 BUFX4_220/Y OAI21X1_466/Y BUFX4_47/Y gnd OAI21X1_467/Y vdd OAI21X1
XOAI21X1_478 INVX2_118/Y BUFX4_164/Y NAND2X1_222/Y gnd OAI21X1_479/B vdd OAI21X1
XOAI21X1_412 NOR2X1_225/Y INVX2_57/Y BUFX4_52/Y gnd AOI21X1_135/C vdd OAI21X1
XOAI21X1_423 BUFX4_221/Y INVX8_19/A INVX1_34/A gnd OAI21X1_427/C vdd OAI21X1
XOAI21X1_445 INVX2_83/Y MUX2X1_6/S OAI21X1_333/C gnd OAI21X1_446/B vdd OAI21X1
XOAI21X1_456 OAI21X1_456/A OAI21X1_456/B OAI21X1_452/Y gnd DFFSR_206/D vdd OAI21X1
XOAI21X1_434 BUFX4_99/Y INVX4_6/Y AND2X2_22/A gnd INVX1_131/A vdd OAI21X1
XOAI21X1_401 BUFX4_222/Y BUFX4_233/Y INVX1_48/A gnd OAI21X1_401/Y vdd OAI21X1
XFILL_35_2_1 gnd vdd FILL
XOAI21X1_83 AND2X2_2/Y INVX1_24/Y NAND3X1_44/Y gnd DFFSR_35/D vdd OAI21X1
XOAI21X1_50 BUFX4_181/Y INVX2_9/Y OAI21X1_50/C gnd DFFSR_1/D vdd OAI21X1
XOAI21X1_61 INVX2_15/Y BUFX4_84/Y OAI21X1_90/C gnd OAI21X1_61/Y vdd OAI21X1
XOAI21X1_72 AND2X2_2/Y INVX1_19/Y OAI21X1_72/C gnd DFFSR_45/D vdd OAI21X1
XOAI21X1_94 INVX2_23/Y BUFX4_11/Y OAI21X1_33/C gnd NAND3X1_51/B vdd OAI21X1
XFILL_26_2_1 gnd vdd FILL
XFILL_1_2_1 gnd vdd FILL
XAND2X2_20 AND2X2_20/A AND2X2_20/B gnd AND2X2_20/Y vdd AND2X2
XOAI21X1_275 OAI21X1_275/A AOI21X1_54/C INVX1_116/A gnd AOI21X1_41/B vdd OAI21X1
XOAI21X1_286 INVX1_104/Y INVX8_13/Y INVX8_9/Y gnd AOI21X1_50/C vdd OAI21X1
XOAI21X1_253 NOR2X1_151/Y NOR2X1_150/Y BUFX4_198/Y gnd OAI21X1_253/Y vdd OAI21X1
XOAI21X1_264 NOR2X1_172/Y NOR2X1_173/Y BUFX4_194/Y gnd OAI21X1_264/Y vdd OAI21X1
XOAI21X1_242 NOR2X1_131/Y NOR2X1_132/Y BUFX4_188/Y gnd OAI21X1_242/Y vdd OAI21X1
XOAI21X1_297 AOI21X1_49/Y AOI21X1_50/Y XOR2X1_4/Y gnd INVX1_125/A vdd OAI21X1
XAND2X2_31 AND2X2_31/A INVX4_9/A gnd AND2X2_31/Y vdd AND2X2
XOAI21X1_220 NOR2X1_99/Y NOR2X1_100/Y AND2X2_15/B gnd OAI21X1_220/Y vdd OAI21X1
XOAI21X1_231 INVX2_165/A BUFX4_238/Y NAND2X1_120/Y gnd AND2X2_16/A vdd OAI21X1
XFILL_9_3_1 gnd vdd FILL
XNAND2X1_270 INVX4_10/A AND2X2_28/A gnd NAND2X1_270/Y vdd NAND2X1
XNAND2X1_281 INVX1_29/A BUFX4_204/Y gnd OAI21X1_647/C vdd NAND2X1
XNAND2X1_292 INVX8_22/A NOR2X1_308/Y gnd NAND2X1_292/Y vdd NAND2X1
XFILL_17_2_1 gnd vdd FILL
XDFFSR_42 DFFSR_42/Q CLKBUF1_27/Y DFFSR_88/R vdd DFFSR_42/D gnd vdd DFFSR
XDFFSR_20 DFFSR_20/Q CLKBUF1_4/Y DFFSR_88/R vdd DFFSR_20/D gnd vdd DFFSR
XDFFSR_64 BUFX2_35/A CLKBUF1_7/Y DFFSR_7/R vdd DFFSR_64/D gnd vdd DFFSR
XDFFSR_53 INVX2_37/A DFFSR_8/CLK DFFSR_53/R vdd DFFSR_53/D gnd vdd DFFSR
XDFFSR_31 INVX1_7/A DFFSR_61/CLK DFFSR_95/R vdd DFFSR_31/D gnd vdd DFFSR
XDFFSR_86 DFFSR_86/Q DFFSR_71/CLK DFFSR_88/R vdd DFFSR_86/D gnd vdd DFFSR
XCLKBUF1_51 CLKBUF1_12/A gnd DFFSR_36/CLK vdd CLKBUF1
XCLKBUF1_40 CLKBUF1_55/Y gnd DFFSR_9/CLK vdd CLKBUF1
XDFFSR_75 BUFX2_46/A DFFSR_59/CLK DFFSR_58/R vdd DFFSR_75/D gnd vdd DFFSR
XDFFSR_97 INVX4_11/A DFFSR_7/CLK DFFSR_98/R vdd DFFSR_97/D gnd vdd DFFSR
XCLKBUF1_62 wb_clk_i gnd CLKBUF1_12/A vdd CLKBUF1
XINVX1_103 INVX1_103/A gnd INVX1_103/Y vdd INVX1
XINVX1_158 INVX1_158/A gnd INVX1_158/Y vdd INVX1
XINVX1_136 INVX1_136/A gnd INVX1_136/Y vdd INVX1
XINVX1_114 INVX1_114/A gnd INVX1_114/Y vdd INVX1
XINVX1_147 INVX1_147/A gnd INVX1_147/Y vdd INVX1
XINVX1_125 INVX1_125/A gnd INVX1_125/Y vdd INVX1
XFILL_32_0_1 gnd vdd FILL
XAOI21X1_118 AOI21X1_118/A AOI21X1_118/B NOR2X1_214/Y gnd DFFSR_231/D vdd AOI21X1
XAOI21X1_107 NOR2X1_207/Y BUFX4_65/Y OAI21X1_337/Y gnd AOI21X1_107/Y vdd AOI21X1
XAOI21X1_129 INVX2_111/Y NAND2X1_234/Y BUFX4_148/Y gnd OAI21X1_394/C vdd AOI21X1
XFILL_23_0_1 gnd vdd FILL
XINVX4_11 INVX4_11/A gnd INVX4_11/Y vdd INVX4
XFILL_6_1_1 gnd vdd FILL
XFILL_14_0_1 gnd vdd FILL
XDFFSR_109 INVX2_41/A CLKBUF1_8/Y vdd BUFX4_89/Y DFFSR_109/D gnd vdd DFFSR
XNOR2X1_324 INVX1_161/A BUFX4_61/Y gnd NOR2X1_324/Y vdd NOR2X1
XNOR2X1_313 INVX1_153/A BUFX4_61/Y gnd NOR2X1_313/Y vdd NOR2X1
XBUFX4_231 BUFX4_230/A gnd BUFX4_231/Y vdd BUFX4
XBUFX4_242 INVX8_16/Y gnd BUFX4_242/Y vdd BUFX4
XNOR2X1_302 BUFX4_30/Y NOR2X1_287/B gnd INVX1_146/A vdd NOR2X1
XBUFX4_220 INVX8_12/Y gnd BUFX4_220/Y vdd BUFX4
XNOR2X1_346 INVX4_5/Y AOI22X1_85/C gnd NOR2X1_346/Y vdd NOR2X1
XFILL_32_2 gnd vdd FILL
XFILL_25_1 gnd vdd FILL
XNOR2X1_335 OR2X2_17/B OR2X2_20/A gnd NOR2X1_335/Y vdd NOR2X1
XNOR2X1_53 NOR2X1_47/Y AND2X2_9/Y gnd INVX2_45/A vdd NOR2X1
XNAND3X1_86 NAND3X1_86/A AOI22X1_1/Y AOI22X1_2/Y gnd DFFSR_81/D vdd NAND3X1
XNAND3X1_42 NAND3X1_42/A BUFX4_15/Y INVX8_2/Y gnd OAI21X1_79/C vdd NAND3X1
XNOR2X1_64 NOR2X1_60/Y NOR2X1_63/Y gnd XOR2X1_2/A vdd NOR2X1
XNAND3X1_64 AND2X2_2/B NAND3X1_64/B BUFX4_107/Y gnd NAND3X1_64/Y vdd NAND3X1
XNAND3X1_31 AND2X2_2/B NAND3X1_31/B BUFX4_27/Y gnd OAI21X1_58/C vdd NAND3X1
XNOR2X1_20 NOR2X1_1/B OAI22X1_4/C gnd INVX8_18/A vdd NOR2X1
XNAND3X1_75 wb_adr_i[3] INVX2_39/Y INVX4_1/Y gnd INVX8_5/A vdd NAND3X1
XNAND3X1_20 BUFX4_20/Y NAND3X1_20/B BUFX4_23/Y gnd OAI21X1_36/C vdd NAND3X1
XNAND3X1_53 BUFX4_20/Y NAND3X1_53/B AND2X2_3/A gnd OAI21X1_99/C vdd NAND3X1
XNOR2X1_42 INVX1_72/Y AND2X2_5/Y gnd NOR2X1_42/Y vdd NOR2X1
XNAND3X1_97 NAND3X1_97/A NAND3X1_97/B NAND3X1_97/C gnd DFFSR_92/D vdd NAND3X1
XNOR2X1_31 NOR3X1_2/A NOR2X1_31/B gnd NOR2X1_31/Y vdd NOR2X1
XNOR2X1_97 INVX2_79/Y NOR2X1_97/B gnd NOR2X1_97/Y vdd NOR2X1
XNOR2X1_86 INVX1_93/Y BUFX4_40/Y gnd NOR2X1_86/Y vdd NOR2X1
XNOR2X1_75 INVX2_61/Y BUFX4_41/Y gnd NOR2X1_75/Y vdd NOR2X1
XNAND2X1_8 MUX2X1_7/S wb_dat_i[31] gnd NAND2X1_8/Y vdd NAND2X1
XNOR2X1_176 NOR2X1_176/A NOR2X1_176/B gnd AOI21X1_36/B vdd NOR2X1
XNOR2X1_154 INVX2_147/Y BUFX4_45/Y gnd NOR2X1_154/Y vdd NOR2X1
XNOR2X1_110 INVX2_93/Y NOR2X1_71/B gnd NOR2X1_110/Y vdd NOR2X1
XNOR2X1_132 INVX2_119/Y BUFX4_46/Y gnd NOR2X1_132/Y vdd NOR2X1
XNOR2X1_143 INVX2_129/Y BUFX4_46/Y gnd NOR2X1_143/Y vdd NOR2X1
XNOR2X1_121 INVX2_110/Y NOR2X1_99/B gnd NOR2X1_121/Y vdd NOR2X1
XNOR2X1_165 INVX2_156/Y BUFX4_41/Y gnd NOR2X1_165/Y vdd NOR2X1
XOAI21X1_649 INVX2_105/Y BUFX4_82/Y OAI21X1_732/C gnd OAI21X1_649/Y vdd OAI21X1
XOAI21X1_605 BUFX4_121/Y OAI21X1_604/Y BUFX4_114/Y gnd OAI21X1_605/Y vdd OAI21X1
XOAI21X1_638 BUFX4_60/Y AOI21X1_237/B OAI21X1_638/C gnd OAI21X1_638/Y vdd OAI21X1
XNOR2X1_198 BUFX4_155/Y AOI21X1_69/C gnd INVX4_10/A vdd NOR2X1
XNOR2X1_187 INVX1_111/Y INVX2_164/Y gnd INVX1_112/A vdd NOR2X1
XOAI21X1_616 AND2X2_30/Y INVX2_85/Y BUFX4_119/Y gnd AOI21X1_219/C vdd OAI21X1
XOAI21X1_627 OAI21X1_627/A OAI21X1_626/Y NAND2X1_275/Y gnd DFFSR_157/D vdd OAI21X1
XINVX1_12 DFFSR_20/Q gnd INVX1_12/Y vdd INVX1
XINVX1_23 INVX2_46/A gnd INVX1_23/Y vdd INVX1
XINVX1_34 INVX1_34/A gnd INVX1_34/Y vdd INVX1
XINVX1_45 INVX1_45/A gnd INVX1_45/Y vdd INVX1
XINVX1_56 INVX1_56/A gnd INVX1_56/Y vdd INVX1
XINVX1_89 INVX1_89/A gnd INVX1_89/Y vdd INVX1
XINVX1_78 INVX1_78/A gnd INVX1_78/Y vdd INVX1
XINVX1_67 INVX2_28/A gnd INVX1_67/Y vdd INVX1
XFILL_31_6_0 gnd vdd FILL
XOAI22X1_18 OAI22X1_9/A INVX1_43/Y INVX8_2/A INVX2_22/Y gnd AOI21X1_7/C vdd OAI22X1
XFILL_22_6_0 gnd vdd FILL
XOAI22X1_29 BUFX4_226/Y INVX1_54/Y INVX8_2/A INVX2_18/Y gnd AOI21X1_12/C vdd OAI22X1
XOAI21X1_413 INVX2_57/Y BUFX4_80/Y NAND2X1_239/Y gnd OAI21X1_414/B vdd OAI21X1
XOAI21X1_468 BUFX4_59/Y AOI21X1_163/B OAI21X1_468/C gnd AOI21X1_164/B vdd OAI21X1
XOAI21X1_479 BUFX4_166/Y OAI21X1_479/B BUFX4_39/Y gnd OAI21X1_480/B vdd OAI21X1
XOAI21X1_424 NOR2X1_228/Y INVX2_114/Y BUFX4_51/Y gnd AOI21X1_140/C vdd OAI21X1
XOAI21X1_435 BUFX4_65/Y NAND2X1_248/Y OAI21X1_435/C gnd AOI21X1_151/B vdd OAI21X1
XOAI21X1_446 BUFX4_168/Y OAI21X1_446/B BUFX4_35/Y gnd OAI21X1_447/B vdd OAI21X1
XOAI21X1_457 BUFX4_67/Y NAND2X1_250/Y AOI21X1_158/Y gnd AOI21X1_159/B vdd OAI21X1
XOAI21X1_402 NOR2X1_223/Y MUX2X1_3/A BUFX4_54/Y gnd AOI21X1_133/C vdd OAI21X1
XFILL_13_6_0 gnd vdd FILL
XOAI21X1_51 INVX2_10/Y BUFX4_82/Y NAND2X1_26/Y gnd NAND3X1_28/B vdd OAI21X1
XOAI21X1_62 BUFX4_181/Y INVX2_15/Y OAI21X1_62/C gnd DFFSR_7/D vdd OAI21X1
XOAI21X1_84 INVX2_19/Y BUFX4_82/Y NAND2X1_28/Y gnd OAI21X1_84/Y vdd OAI21X1
XOAI21X1_40 BUFX4_182/Y INVX2_4/Y OAI21X1_40/C gnd DFFSR_12/D vdd OAI21X1
XOAI21X1_73 BUFX4_91/Y BUFX4_9/Y OAI21X1_73/C gnd OAI21X1_73/Y vdd OAI21X1
XOAI21X1_95 AND2X2_3/Y INVX2_23/Y OAI21X1_95/C gnd DFFSR_55/D vdd OAI21X1
XOAI21X1_210 NOR2X1_80/Y NOR2X1_79/Y BUFX4_195/Y gnd OAI21X1_210/Y vdd OAI21X1
XOAI21X1_221 NOR2X1_101/Y NOR2X1_102/Y BUFX4_197/Y gnd OAI21X1_221/Y vdd OAI21X1
XOAI21X1_276 INVX2_51/Y INVX8_13/Y INVX8_9/Y gnd AOI21X1_42/C vdd OAI21X1
XAND2X2_10 AND2X2_10/A NOR2X1_58/Y gnd AND2X2_10/Y vdd AND2X2
XAND2X2_21 AND2X2_21/A AND2X2_21/B gnd AND2X2_21/Y vdd AND2X2
XOAI21X1_287 INVX1_89/Y INVX1_17/A AOI21X1_32/Y gnd OAI21X1_287/Y vdd OAI21X1
XOAI21X1_254 NOR2X1_153/Y NOR2X1_152/Y BUFX4_184/Y gnd NAND3X1_156/C vdd OAI21X1
XOAI21X1_265 OR2X2_3/B NOR2X1_51/A BUFX2_1/A gnd NAND2X1_127/A vdd OAI21X1
XAND2X2_32 AND2X2_32/A INVX4_8/A gnd AND2X2_32/Y vdd AND2X2
XOAI21X1_298 INVX4_11/A INVX1_17/A NAND2X1_170/Y gnd AOI21X1_68/C vdd OAI21X1
XOAI21X1_243 NOR2X1_133/Y NOR2X1_134/Y BUFX4_197/Y gnd OAI21X1_243/Y vdd OAI21X1
XOAI21X1_232 AND2X2_15/Y AND2X2_16/Y BUFX4_41/Y gnd OAI21X1_232/Y vdd OAI21X1
XNAND2X1_282 INVX1_27/A BUFX4_204/Y gnd OAI21X1_651/C vdd NAND2X1
XNAND2X1_293 INVX2_161/Y NAND2X1_292/Y gnd NAND2X1_293/Y vdd NAND2X1
XNAND2X1_260 INVX2_109/A BUFX4_207/Y gnd NAND2X1_260/Y vdd NAND2X1
XNAND2X1_271 INVX4_10/A NOR2X1_266/Y gnd AOI21X1_216/B vdd NAND2X1
XDFFSR_65 DFFSR_65/Q CLKBUF1_4/Y DFFSR_88/R vdd DFFSR_65/D gnd vdd DFFSR
XDFFSR_21 INVX1_13/A DFFSR_6/CLK DFFSR_1/R vdd DFFSR_21/D gnd vdd DFFSR
XDFFSR_87 BUFX2_58/A DFFSR_87/CLK DFFSR_9/R vdd DFFSR_87/D gnd vdd DFFSR
XDFFSR_54 DFFSR_54/Q DFFSR_9/CLK DFFSR_9/R vdd DFFSR_54/D gnd vdd DFFSR
XDFFSR_43 DFFSR_43/Q CLKBUF1_23/Y DFFSR_53/R vdd DFFSR_43/D gnd vdd DFFSR
XDFFSR_10 INVX2_2/A CLKBUF1_35/Y DFFSR_53/R vdd DFFSR_10/D gnd vdd DFFSR
XDFFSR_76 BUFX2_47/A DFFSR_46/CLK DFFSR_58/R vdd DFFSR_76/D gnd vdd DFFSR
XDFFSR_32 INVX1_8/A DFFSR_47/CLK DFFSR_95/R vdd DFFSR_32/D gnd vdd DFFSR
XDFFSR_98 DFFSR_98/Q DFFSR_98/CLK DFFSR_98/R vdd DFFSR_98/D gnd vdd DFFSR
XCLKBUF1_41 CLKBUF1_7/A gnd DFFSR_8/CLK vdd CLKBUF1
XCLKBUF1_30 CLKBUF1_34/A gnd DFFSR_26/CLK vdd CLKBUF1
XCLKBUF1_52 CLKBUF1_34/A gnd CLKBUF1_52/Y vdd CLKBUF1
XCLKBUF1_63 wb_clk_i gnd DFFSR_59/CLK vdd CLKBUF1
XFILL_27_5_0 gnd vdd FILL
XFILL_2_5_0 gnd vdd FILL
XFILL_10_4_0 gnd vdd FILL
XINVX1_115 INVX1_115/A gnd INVX1_115/Y vdd INVX1
XINVX1_104 OR2X2_8/B gnd INVX1_104/Y vdd INVX1
XINVX1_159 INVX1_159/A gnd INVX1_159/Y vdd INVX1
XINVX1_137 INVX1_137/A gnd INVX1_137/Y vdd INVX1
XINVX1_148 INVX1_148/A gnd INVX1_148/Y vdd INVX1
XINVX1_126 INVX1_126/A gnd INVX1_126/Y vdd INVX1
XFILL_18_5_0 gnd vdd FILL
XAOI21X1_119 NOR2X1_215/Y BUFX4_59/Y AOI21X1_119/C gnd OAI21X1_374/A vdd AOI21X1
XAOI21X1_108 NOR2X1_208/Y BUFX4_65/Y AOI21X1_108/C gnd OAI21X1_345/A vdd AOI21X1
XNOR2X1_347 NOR2X1_347/A NOR2X1_347/B gnd AOI22X1_85/A vdd NOR2X1
XFILL_32_3 gnd vdd FILL
XNOR2X1_336 INVX1_44/A BUFX4_244/Y gnd NOR2X1_336/Y vdd NOR2X1
XBUFX4_232 BUFX4_230/A gnd INVX8_19/A vdd BUFX4
XNOR2X1_314 OR2X2_18/B NOR2X1_296/B gnd INVX1_154/A vdd NOR2X1
XNOR2X1_325 INVX4_7/Y NOR2X1_329/B gnd NOR2X1_325/Y vdd NOR2X1
XBUFX4_210 BUFX4_211/A gnd BUFX4_210/Y vdd BUFX4
XNOR2X1_303 INVX8_22/Y INVX1_146/Y gnd INVX1_147/A vdd NOR2X1
XBUFX4_243 INVX8_16/Y gnd BUFX4_243/Y vdd BUFX4
XBUFX4_221 INVX8_12/Y gnd BUFX4_221/Y vdd BUFX4
XFILL_33_3_0 gnd vdd FILL
XFILL_25_2 gnd vdd FILL
XFILL_24_3_0 gnd vdd FILL
XNAND3X1_32 BUFX4_16/Y OAI21X1_59/Y BUFX4_24/Y gnd OAI21X1_60/C vdd NAND3X1
XNAND3X1_10 BUFX4_14/Y NAND3X1_10/B BUFX4_23/Y gnd OAI21X1_16/C vdd NAND3X1
XFILL_7_4_0 gnd vdd FILL
XNAND3X1_21 AND2X2_1/B NAND3X1_21/B BUFX4_23/Y gnd OAI21X1_38/C vdd NAND3X1
XNOR2X1_65 OR2X2_7/B INVX2_50/Y gnd NOR2X1_65/Y vdd NOR2X1
XNAND3X1_87 NAND3X1_87/A AOI22X1_3/Y AOI22X1_4/Y gnd DFFSR_82/D vdd NAND3X1
XNAND3X1_43 NAND3X1_43/A BUFX4_15/Y INVX8_2/Y gnd OAI21X1_81/C vdd NAND3X1
XNOR2X1_54 XNOR2X1_3/Y INVX1_81/Y gnd NOR2X1_54/Y vdd NOR2X1
XNOR2X1_10 NOR2X1_10/A NOR2X1_10/B gnd NOR2X1_10/Y vdd NOR2X1
XNAND3X1_65 BUFX4_18/Y NAND3X1_65/B BUFX4_106/Y gnd NAND3X1_65/Y vdd NAND3X1
XNAND3X1_76 wb_adr_i[3] INVX2_134/A NOR2X1_4/Y gnd NAND2X1_46/A vdd NAND3X1
XNAND3X1_54 AND2X2_1/B NAND3X1_54/B BUFX4_108/Y gnd NAND3X1_54/Y vdd NAND3X1
XNAND3X1_98 NAND3X1_98/A NAND3X1_98/B NAND3X1_98/C gnd DFFSR_93/D vdd NAND3X1
XNOR2X1_43 INVX1_74/Y NOR2X1_40/Y gnd NOR2X1_43/Y vdd NOR2X1
XNOR2X1_87 INVX2_70/Y NOR2X1_87/B gnd NOR2X1_87/Y vdd NOR2X1
XNOR2X1_32 INVX2_29/A INVX2_30/A gnd NOR2X1_32/Y vdd NOR2X1
XNOR2X1_21 NOR2X1_1/B INVX8_5/A gnd INVX8_11/A vdd NOR2X1
XNOR2X1_76 INVX2_62/Y NOR2X1_76/B gnd NOR2X1_76/Y vdd NOR2X1
XNOR2X1_98 INVX2_80/Y BUFX4_44/Y gnd NOR2X1_98/Y vdd NOR2X1
XFILL_15_3_0 gnd vdd FILL
XNAND2X1_9 wb_dat_i[16] NAND2X1_9/B gnd NAND2X1_9/Y vdd NAND2X1
XNOR2X1_177 INVX2_42/A NOR2X1_177/B gnd NOR2X1_177/Y vdd NOR2X1
XNOR2X1_155 INVX2_148/Y BUFX4_217/Y gnd NOR2X1_155/Y vdd NOR2X1
XNOR2X1_166 INVX2_157/Y NOR2X1_97/B gnd NOR2X1_166/Y vdd NOR2X1
XNOR2X1_111 INVX2_94/Y BUFX4_42/Y gnd NOR2X1_111/Y vdd NOR2X1
XNOR2X1_144 INVX2_130/Y BUFX4_215/Y gnd NOR2X1_144/Y vdd NOR2X1
XNOR2X1_133 INVX2_120/Y BUFX4_215/Y gnd NOR2X1_133/Y vdd NOR2X1
XNOR2X1_199 XOR2X1_4/Y INVX1_110/Y gnd INVX1_122/A vdd NOR2X1
XNOR2X1_122 INVX1_96/Y BUFX4_43/Y gnd NOR2X1_122/Y vdd NOR2X1
XNOR2X1_188 INVX8_14/Y INVX1_112/Y gnd NOR2X1_188/Y vdd NOR2X1
XNOR2X1_100 INVX1_95/Y BUFX4_43/Y gnd NOR2X1_100/Y vdd NOR2X1
XOAI21X1_606 OAI21X1_606/A OAI21X1_605/Y OAI21X1_606/C gnd DFFSR_165/D vdd OAI21X1
XOAI21X1_639 INVX2_115/Y BUFX4_79/Y NAND2X1_243/Y gnd AOI21X1_238/B vdd OAI21X1
XOAI21X1_628 BUFX4_64/Y OAI21X1_628/B AOI21X1_227/Y gnd OAI21X1_628/Y vdd OAI21X1
XOAI21X1_617 INVX2_85/Y BUFX4_10/Y OAI21X1_699/C gnd OAI21X1_618/B vdd OAI21X1
XINVX1_13 INVX1_13/A gnd INVX1_13/Y vdd INVX1
XINVX1_24 INVX4_2/A gnd INVX1_24/Y vdd INVX1
XINVX1_79 INVX1_79/A gnd INVX1_79/Y vdd INVX1
XINVX1_35 INVX1_35/A gnd INVX1_35/Y vdd INVX1
XINVX1_46 INVX1_46/A gnd INVX1_46/Y vdd INVX1
XINVX1_57 INVX1_57/A gnd INVX1_57/Y vdd INVX1
XINVX1_68 DFFSR_57/Q gnd INVX1_68/Y vdd INVX1
XFILL_31_6_1 gnd vdd FILL
XFILL_30_1_0 gnd vdd FILL
XFILL_22_6_1 gnd vdd FILL
XOAI22X1_19 INVX8_1/A INVX2_16/Y INVX1_44/Y OAI22X1_9/A gnd NOR2X1_11/A vdd OAI22X1
XFILL_21_1_0 gnd vdd FILL
XOAI21X1_414 BUFX4_52/Y OAI21X1_414/B BUFX4_244/Y gnd OAI21X1_415/B vdd OAI21X1
XOAI21X1_403 MUX2X1_3/A BUFX4_6/Y OAI21X1_515/C gnd OAI21X1_404/B vdd OAI21X1
XOAI21X1_425 INVX2_114/Y BUFX4_86/Y NAND2X1_243/Y gnd OAI21X1_426/B vdd OAI21X1
XOAI21X1_469 INVX2_160/Y BUFX4_162/Y NAND2X1_216/Y gnd OAI21X1_470/B vdd OAI21X1
XOAI21X1_436 INVX2_66/Y BUFX4_72/Y OAI21X1_323/C gnd OAI21X1_437/B vdd OAI21X1
XOAI21X1_447 OAI21X1_447/A OAI21X1_447/B OAI21X1_442/Y gnd DFFSR_208/D vdd OAI21X1
XOAI21X1_458 MUX2X1_4/B BUFX4_70/Y OAI21X1_458/C gnd OAI21X1_458/Y vdd OAI21X1
XFILL_29_2_0 gnd vdd FILL
XFILL_4_2_0 gnd vdd FILL
XFILL_12_1_0 gnd vdd FILL
XFILL_13_6_1 gnd vdd FILL
XOAI21X1_52 BUFX4_181/Y INVX2_10/Y NAND3X1_28/Y gnd DFFSR_2/D vdd OAI21X1
XOAI21X1_30 BUFX4_179/Y INVX1_15/Y OAI21X1_30/C gnd DFFSR_23/D vdd OAI21X1
XOAI21X1_63 INVX2_16/Y BUFX4_86/Y OAI21X1_92/C gnd NAND3X1_34/B vdd OAI21X1
XOAI21X1_41 INVX2_5/Y BUFX4_6/Y OAI21X1_71/C gnd NAND3X1_23/B vdd OAI21X1
XOAI21X1_85 AND2X2_2/Y INVX2_19/Y NAND3X1_45/Y gnd DFFSR_36/D vdd OAI21X1
XOAI21X1_74 AND2X2_2/Y BUFX4_91/Y OAI21X1_74/C gnd DFFSR_46/D vdd OAI21X1
XOAI21X1_96 INVX2_24/Y BUFX4_12/Y OAI21X1_65/C gnd NAND3X1_52/B vdd OAI21X1
XOAI21X1_255 NOR2X1_155/Y NOR2X1_154/Y BUFX4_198/Y gnd NAND3X1_157/B vdd OAI21X1
XOAI21X1_233 NOR2X1_113/Y NOR2X1_114/Y BUFX4_198/Y gnd OAI21X1_233/Y vdd OAI21X1
XOAI21X1_200 AND2X2_11/A NAND2X1_110/Y AOI21X1_29/Y gnd OR2X2_9/A vdd OAI21X1
XOAI21X1_211 NOR2X1_82/Y NOR2X1_81/Y AND2X2_15/B gnd OAI21X1_211/Y vdd OAI21X1
XOAI21X1_244 NOR2X1_135/Y NOR2X1_136/Y AND2X2_16/B gnd NAND3X1_148/B vdd OAI21X1
XOAI21X1_222 NOR2X1_103/Y NOR2X1_104/Y BUFX4_188/Y gnd OAI21X1_222/Y vdd OAI21X1
XAND2X2_33 AND2X2_33/A AND2X2_33/B gnd AND2X2_33/Y vdd AND2X2
XOAI21X1_288 AOI21X1_51/Y INVX1_105/A BUFX4_248/Y gnd OAI21X1_289/A vdd OAI21X1
XAND2X2_11 AND2X2_11/A INVX1_87/Y gnd AND2X2_11/Y vdd AND2X2
XOAI21X1_277 AOI21X1_44/Y NOR2X1_181/Y OAI21X1_277/C gnd OAI21X1_277/Y vdd OAI21X1
XOAI21X1_266 INVX8_18/A NOR2X1_19/Y INVX4_5/Y gnd BUFX4_36/A vdd OAI21X1
XAND2X2_22 AND2X2_22/A INVX8_14/A gnd AND2X2_22/Y vdd AND2X2
XOAI21X1_299 INVX2_86/A BUFX4_175/Y AOI21X1_73/Y gnd NAND3X1_202/A vdd OAI21X1
XNAND2X1_294 BUFX4_204/Y OAI21X1_672/Y gnd NAND2X1_294/Y vdd NAND2X1
XNAND2X1_283 BUFX4_207/Y NAND2X1_283/B gnd OAI21X1_655/C vdd NAND2X1
XNAND2X1_261 INVX2_68/A BUFX4_205/Y gnd NAND2X1_261/Y vdd NAND2X1
XNAND2X1_250 INVX4_7/A AND2X2_24/A gnd NAND2X1_250/Y vdd NAND2X1
XNAND2X1_272 INVX1_56/A BUFX4_203/Y gnd NAND2X1_272/Y vdd NAND2X1
XFILL_6_1 gnd vdd FILL
XFILL_35_0_0 gnd vdd FILL
XDFFSR_88 DFFSR_88/Q DFFSR_88/CLK DFFSR_88/R vdd DFFSR_88/D gnd vdd DFFSR
XDFFSR_22 DFFSR_22/Q DFFSR_82/CLK DFFSR_2/R vdd DFFSR_22/D gnd vdd DFFSR
XDFFSR_77 BUFX2_48/A DFFSR_2/CLK DFFSR_7/R vdd DFFSR_77/D gnd vdd DFFSR
XDFFSR_66 BUFX2_37/A DFFSR_6/CLK DFFSR_7/R vdd DFFSR_66/D gnd vdd DFFSR
XDFFSR_33 DFFSR_33/Q DFFSR_3/CLK DFFSR_7/R vdd DFFSR_33/D gnd vdd DFFSR
XDFFSR_44 DFFSR_44/Q CLKBUF1_5/A DFFSR_53/R vdd DFFSR_44/D gnd vdd DFFSR
XDFFSR_55 DFFSR_55/Q CLKBUF1_35/Y DFFSR_58/R vdd DFFSR_55/D gnd vdd DFFSR
XDFFSR_11 INVX2_3/A DFFSR_56/CLK DFFSR_95/R vdd DFFSR_11/D gnd vdd DFFSR
XDFFSR_99 BUFX2_2/A DFFSR_99/CLK DFFSR_98/R vdd DFFSR_99/D gnd vdd DFFSR
XCLKBUF1_53 wb_clk_i gnd CLKBUF1_46/A vdd CLKBUF1
XCLKBUF1_64 wb_clk_i gnd CLKBUF1_7/A vdd CLKBUF1
XCLKBUF1_20 CLKBUF1_38/A gnd DFFSR_61/CLK vdd CLKBUF1
XCLKBUF1_42 CLKBUF1_34/A gnd CLKBUF1_42/Y vdd CLKBUF1
XCLKBUF1_31 CLKBUF1_5/A gnd DFFSR_56/CLK vdd CLKBUF1
XFILL_27_5_1 gnd vdd FILL
XFILL_26_0_0 gnd vdd FILL
XFILL_2_5_1 gnd vdd FILL
XFILL_1_0_0 gnd vdd FILL
XINVX1_116 INVX1_116/A gnd INVX1_116/Y vdd INVX1
XINVX1_105 INVX1_105/A gnd INVX1_105/Y vdd INVX1
XFILL_10_4_1 gnd vdd FILL
XINVX1_149 INVX1_149/A gnd INVX1_149/Y vdd INVX1
XINVX1_127 INVX1_127/A gnd INVX1_127/Y vdd INVX1
XINVX1_138 DFFSR_172/Q gnd INVX1_138/Y vdd INVX1
XFILL_9_1_0 gnd vdd FILL
XFILL_18_5_1 gnd vdd FILL
XFILL_17_0_0 gnd vdd FILL
XAOI21X1_109 NOR2X1_209/Y BUFX4_65/Y AOI21X1_109/C gnd OAI21X1_350/A vdd AOI21X1
XBUFX4_211 BUFX4_211/A gnd BUFX4_211/Y vdd BUFX4
XBUFX4_200 BUFX4_200/A gnd OAI22X1_4/A vdd BUFX4
XNOR2X1_348 INVX2_46/A DFFSR_33/Q gnd AND2X2_33/B vdd NOR2X1
XFILL_33_3_1 gnd vdd FILL
XFILL_25_3 gnd vdd FILL
XBUFX4_244 INVX8_16/Y gnd BUFX4_244/Y vdd BUFX4
XNOR2X1_304 INVX1_147/Y BUFX4_63/Y gnd NOR2X1_304/Y vdd NOR2X1
XNOR2X1_337 OR2X2_18/B NOR2X1_337/B gnd INVX1_163/A vdd NOR2X1
XNOR2X1_326 OR2X2_12/A INVX1_112/Y gnd NOR2X1_326/Y vdd NOR2X1
XNOR2X1_315 INVX1_154/Y BUFX4_62/Y gnd NOR2X1_315/Y vdd NOR2X1
XBUFX4_222 INVX8_12/Y gnd BUFX4_222/Y vdd BUFX4
XBUFX4_233 BUFX4_230/A gnd BUFX4_233/Y vdd BUFX4
XFILL_24_3_1 gnd vdd FILL
XNAND3X1_11 BUFX4_19/Y NAND3X1_11/B BUFX4_26/Y gnd OAI21X1_18/C vdd NAND3X1
XNAND3X1_44 NAND3X1_44/A BUFX4_16/Y INVX8_2/Y gnd NAND3X1_44/Y vdd NAND3X1
XNAND3X1_33 BUFX4_15/Y OAI21X1_61/Y BUFX4_24/Y gnd OAI21X1_62/C vdd NAND3X1
XNAND3X1_66 AND2X2_2/B NAND3X1_66/B BUFX4_106/Y gnd NAND3X1_66/Y vdd NAND3X1
XNAND3X1_22 BUFX4_20/Y OAI21X1_39/Y BUFX4_23/Y gnd OAI21X1_40/C vdd NAND3X1
XNAND3X1_55 AND2X2_1/B NAND3X1_55/B AND2X2_3/A gnd NAND3X1_55/Y vdd NAND3X1
XFILL_7_4_1 gnd vdd FILL
XNOR2X1_66 INVX2_50/A INVX2_51/Y gnd NOR2X1_67/B vdd NOR2X1
XNOR2X1_55 XNOR2X1_4/Y NOR2X1_55/B gnd NOR2X1_55/Y vdd NOR2X1
XNAND3X1_88 AOI22X1_6/Y NAND2X1_62/Y AOI22X1_5/Y gnd DFFSR_83/D vdd NAND3X1
XNAND3X1_77 wb_adr_i[4] DFFSR_40/Q NOR2X1_3/Y gnd NAND2X1_46/B vdd NAND3X1
XNOR2X1_11 NOR2X1_11/A NOR2X1_11/B gnd NOR2X1_11/Y vdd NOR2X1
XNOR2X1_22 NOR2X1_1/B OAI22X1_9/A gnd INVX4_6/A vdd NOR2X1
XFILL_15_3_1 gnd vdd FILL
XNAND3X1_99 NAND3X1_99/A NAND3X1_99/B NAND3X1_99/C gnd DFFSR_94/D vdd NAND3X1
XNOR2X1_99 INVX2_83/Y NOR2X1_99/B gnd NOR2X1_99/Y vdd NOR2X1
XNOR2X1_44 OR2X2_4/A NOR2X1_44/B gnd NOR2X1_44/Y vdd NOR2X1
XNOR2X1_88 INVX2_71/Y BUFX4_40/Y gnd NOR2X1_88/Y vdd NOR2X1
XNOR2X1_77 INVX1_91/Y BUFX4_41/Y gnd NOR2X1_77/Y vdd NOR2X1
XNOR2X1_33 DFFSR_55/Q INVX2_24/A gnd NOR2X1_33/Y vdd NOR2X1
XNOR2X1_178 INVX2_49/Y OR2X2_11/A gnd NOR2X1_178/Y vdd NOR2X1
XNOR2X1_156 INVX1_100/Y BUFX4_45/Y gnd NOR2X1_156/Y vdd NOR2X1
XNOR2X1_167 INVX1_102/Y BUFX4_44/Y gnd NOR2X1_167/Y vdd NOR2X1
XNOR2X1_112 INVX2_95/Y NOR2X1_71/B gnd NOR2X1_112/Y vdd NOR2X1
XNOR2X1_189 INVX1_114/Y INVX1_113/Y gnd NOR2X1_189/Y vdd NOR2X1
XNOR2X1_145 INVX2_131/Y BUFX4_46/Y gnd NOR2X1_145/Y vdd NOR2X1
XNOR2X1_134 INVX2_121/Y BUFX4_46/Y gnd NOR2X1_134/Y vdd NOR2X1
XNOR2X1_123 INVX2_111/Y NOR2X1_87/B gnd NOR2X1_123/Y vdd NOR2X1
XNOR2X1_101 INVX2_84/Y BUFX4_215/Y gnd NOR2X1_101/Y vdd NOR2X1
XOAI21X1_607 BUFX4_98/Y INVX8_11/Y AND2X2_27/A gnd NOR2X1_282/B vdd OAI21X1
XOAI21X1_618 BUFX4_120/Y OAI21X1_618/B BUFX4_118/Y gnd OAI21X1_619/B vdd OAI21X1
XOAI21X1_629 INVX2_97/Y BUFX4_6/Y NAND2X1_238/Y gnd AOI21X1_228/B vdd OAI21X1
XINVX1_14 DFFSR_22/Q gnd INVX1_14/Y vdd INVX1
XINVX1_25 DFFSR_40/Q gnd INVX1_25/Y vdd INVX1
XINVX1_36 INVX1_36/A gnd INVX1_36/Y vdd INVX1
XINVX1_47 INVX1_47/A gnd INVX1_47/Y vdd INVX1
XINVX1_58 INVX1_58/A gnd INVX1_58/Y vdd INVX1
XINVX1_69 INVX2_26/A gnd INVX1_69/Y vdd INVX1
XFILL_30_1_1 gnd vdd FILL
XFILL_21_1_1 gnd vdd FILL
XOAI21X1_426 BUFX4_52/Y OAI21X1_426/B BUFX4_244/Y gnd OAI21X1_427/B vdd OAI21X1
XOAI21X1_415 OAI21X1_415/A OAI21X1_415/B OAI21X1_411/Y gnd DFFSR_218/D vdd OAI21X1
XOAI21X1_437 BUFX4_223/Y OAI21X1_437/B BUFX4_50/Y gnd AOI21X1_151/A vdd OAI21X1
XOAI21X1_448 BUFX4_99/Y INVX4_6/Y INVX1_130/Y gnd INVX1_133/A vdd OAI21X1
XOAI21X1_404 BUFX4_54/Y OAI21X1_404/B BUFX4_243/Y gnd OAI21X1_405/B vdd OAI21X1
XDFFSR_250 INVX2_42/A DFFSR_85/CLK DFFSR_165/R vdd DFFSR_250/D gnd vdd DFFSR
XOAI21X1_459 BUFX4_224/Y OAI21X1_458/Y BUFX4_50/Y gnd AOI21X1_159/A vdd OAI21X1
XFILL_29_2_1 gnd vdd FILL
XFILL_4_2_1 gnd vdd FILL
XFILL_12_1_1 gnd vdd FILL
XINVX2_90 INVX2_90/A gnd INVX2_90/Y vdd INVX2
XOAI21X1_31 INVX1_16/Y BUFX4_160/Y OAI21X1_31/C gnd NAND3X1_18/B vdd OAI21X1
XOAI21X1_20 BUFX4_181/Y INVX1_10/Y NAND3X1_12/Y gnd DFFSR_18/D vdd OAI21X1
XOAI21X1_53 INVX2_11/Y BUFX4_84/Y NAND2X1_27/Y gnd OAI21X1_53/Y vdd OAI21X1
XOAI21X1_86 INVX2_20/Y BUFX4_83/Y OAI21X1_86/C gnd NAND3X1_46/A vdd OAI21X1
XOAI21X1_64 BUFX4_183/Y INVX2_16/Y OAI21X1_64/C gnd DFFSR_8/D vdd OAI21X1
XOAI21X1_75 INVX1_20/Y BUFX4_10/Y OAI21X1_33/C gnd OAI21X1_75/Y vdd OAI21X1
XOAI21X1_42 BUFX4_183/Y INVX2_5/Y OAI21X1_42/C gnd DFFSR_13/D vdd OAI21X1
XOAI21X1_97 AND2X2_3/Y INVX2_24/Y OAI21X1_97/C gnd DFFSR_56/D vdd OAI21X1
XOAI21X1_278 AOI21X1_45/Y NOR2X1_178/Y AOI21X1_37/C gnd NAND3X1_191/C vdd OAI21X1
XOAI21X1_289 OAI21X1_289/A INVX1_115/Y OAI21X1_287/Y gnd BUFX4_154/A vdd OAI21X1
XOAI21X1_256 NOR2X1_157/Y NOR2X1_156/Y BUFX4_184/Y gnd NAND3X1_157/C vdd OAI21X1
XOAI21X1_201 AND2X2_12/Y NOR2X1_68/Y INVX8_9/A gnd OAI21X1_202/C vdd OAI21X1
XOAI21X1_234 NOR2X1_115/Y NOR2X1_116/Y BUFX4_198/Y gnd OAI21X1_234/Y vdd OAI21X1
XOAI21X1_223 NOR2X1_106/Y NOR2X1_105/Y BUFX4_197/Y gnd NAND3X1_129/B vdd OAI21X1
XOAI21X1_267 BUFX4_224/Y BUFX4_231/Y DFFSR_243/Q gnd OAI21X1_267/Y vdd OAI21X1
XOAI21X1_212 NOR2X1_83/Y NOR2X1_84/Y BUFX4_195/Y gnd OAI21X1_212/Y vdd OAI21X1
XOAI21X1_245 NOR2X1_137/Y NOR2X1_138/Y BUFX4_187/Y gnd OAI21X1_245/Y vdd OAI21X1
XAND2X2_12 OR2X2_9/A OR2X2_9/B gnd AND2X2_12/Y vdd AND2X2
XAND2X2_23 AND2X2_23/A INVX4_7/A gnd AND2X2_23/Y vdd AND2X2
XNAND2X1_240 BUFX4_81/Y wb_dat_i[5] gnd NAND2X1_240/Y vdd NAND2X1
XNAND2X1_251 INVX4_7/A AND2X2_25/A gnd OAI21X1_465/B vdd NAND2X1
XNAND2X1_295 INVX8_21/A NAND2X1_295/B gnd OAI21X1_678/C vdd NAND2X1
XNAND2X1_262 DFFSR_173/Q BUFX4_207/Y gnd NAND2X1_262/Y vdd NAND2X1
XNAND2X1_284 INVX1_142/A BUFX4_62/Y gnd AOI22X1_78/C vdd NAND2X1
XNAND2X1_273 INVX4_10/A AND2X2_29/A gnd AOI21X1_220/B vdd NAND2X1
XOAI21X1_790 OAI21X1_790/A BUFX4_206/Y NAND2X1_340/Y gnd DFFSR_123/D vdd OAI21X1
XFILL_35_0_1 gnd vdd FILL
XDFFSR_12 INVX2_4/A DFFSR_87/CLK DFFSR_53/R vdd DFFSR_12/D gnd vdd DFFSR
XDFFSR_67 BUFX2_38/A DFFSR_82/CLK DFFSR_2/R vdd DFFSR_67/D gnd vdd DFFSR
XDFFSR_23 INVX1_15/A DFFSR_83/CLK DFFSR_1/R vdd DFFSR_23/D gnd vdd DFFSR
XDFFSR_34 INVX2_46/A CLKBUF1_7/Y DFFSR_7/R vdd DFFSR_34/D gnd vdd DFFSR
XDFFSR_45 INVX1_19/A CLKBUF1_5/A DFFSR_53/R vdd DFFSR_45/D gnd vdd DFFSR
XDFFSR_78 BUFX2_49/A DFFSR_78/CLK DFFSR_58/R vdd DFFSR_78/D gnd vdd DFFSR
XDFFSR_89 DFFSR_89/Q CLKBUF1_34/A DFFSR_25/R vdd DFFSR_89/D gnd vdd DFFSR
XDFFSR_56 INVX2_24/A DFFSR_56/CLK DFFSR_58/R vdd DFFSR_56/D gnd vdd DFFSR
XCLKBUF1_54 wb_clk_i gnd CLKBUF1_54/Y vdd CLKBUF1
XCLKBUF1_65 wb_clk_i gnd CLKBUF1_6/A vdd CLKBUF1
XCLKBUF1_32 CLKBUF1_32/A gnd CLKBUF1_32/Y vdd CLKBUF1
XCLKBUF1_10 CLKBUF1_38/A gnd DFFSR_78/CLK vdd CLKBUF1
XCLKBUF1_43 CLKBUF1_5/A gnd DFFSR_98/CLK vdd CLKBUF1
XCLKBUF1_21 DFFSR_59/CLK gnd DFFSR_28/CLK vdd CLKBUF1
XFILL_26_0_1 gnd vdd FILL
XFILL_1_0_1 gnd vdd FILL
XINVX1_106 INVX1_106/A gnd INVX1_106/Y vdd INVX1
XINVX1_117 INVX1_117/A gnd INVX1_117/Y vdd INVX1
XINVX1_128 INVX1_128/A gnd INVX1_128/Y vdd INVX1
XINVX1_139 INVX1_139/A gnd INVX1_139/Y vdd INVX1
XFILL_9_1_1 gnd vdd FILL
XFILL_17_0_1 gnd vdd FILL
XBUFX4_245 DFFSR_44/Q gnd BUFX4_245/Y vdd BUFX4
XBUFX4_201 BUFX4_200/A gnd OAI22X1_7/D vdd BUFX4
XBUFX4_223 INVX8_12/Y gnd BUFX4_223/Y vdd BUFX4
XBUFX4_234 BUFX4_230/A gnd BUFX4_234/Y vdd BUFX4
XBUFX4_212 BUFX4_211/A gnd BUFX4_212/Y vdd BUFX4
XNOR2X1_349 NOR2X1_50/A INVX4_5/Y gnd AOI22X1_85/D vdd NOR2X1
XNOR2X1_327 OR2X2_21/B INVX8_14/Y gnd NOR2X1_327/Y vdd NOR2X1
XNOR2X1_305 INVX8_22/Y OR2X2_19/A gnd INVX1_148/A vdd NOR2X1
XNOR2X1_338 INVX1_163/Y BUFX4_63/Y gnd NOR2X1_338/Y vdd NOR2X1
XNOR2X1_316 OR2X2_18/B NOR2X1_316/B gnd INVX1_155/A vdd NOR2X1
XNAND3X1_12 BUFX4_16/Y NAND3X1_12/B BUFX4_24/Y gnd NAND3X1_12/Y vdd NAND3X1
XNAND3X1_45 OAI21X1_84/Y BUFX4_16/Y INVX8_2/Y gnd NAND3X1_45/Y vdd NAND3X1
XNAND3X1_34 AND2X2_2/B NAND3X1_34/B BUFX4_27/Y gnd OAI21X1_64/C vdd NAND3X1
XNAND3X1_67 wb_adr_i[2] wb_adr_i[3] INVX2_39/Y gnd BUFX4_228/A vdd NAND3X1
XNAND3X1_89 NAND2X1_63/Y AOI22X1_7/Y AOI22X1_8/Y gnd DFFSR_84/D vdd NAND3X1
XNAND3X1_23 BUFX4_20/Y NAND3X1_23/B BUFX4_27/Y gnd OAI21X1_42/C vdd NAND3X1
XNOR2X1_12 NOR2X1_12/A NOR2X1_12/B gnd NOR2X1_12/Y vdd NOR2X1
XNAND3X1_56 BUFX4_20/Y NAND3X1_56/B AND2X2_3/A gnd NAND3X1_56/Y vdd NAND3X1
XNAND3X1_78 wb_adr_i[3] INVX2_98/A NOR2X1_4/Y gnd NAND3X1_78/Y vdd NAND3X1
XNOR2X1_56 INVX2_48/A INVX4_3/Y gnd NOR2X1_56/Y vdd NOR2X1
XNOR2X1_67 NOR2X1_65/Y NOR2X1_67/B gnd XOR2X1_2/B vdd NOR2X1
XNOR2X1_23 INVX2_41/A INVX1_75/A gnd AND2X2_8/B vdd NOR2X1
XNOR2X1_45 NOR2X1_44/Y BUFX4_2/Y gnd NOR2X1_45/Y vdd NOR2X1
XNOR2X1_89 INVX2_72/Y NOR2X1_76/B gnd NOR2X1_89/Y vdd NOR2X1
XNOR2X1_78 INVX2_63/Y NOR2X1_76/B gnd NOR2X1_78/Y vdd NOR2X1
XNOR2X1_34 NOR2X1_34/A NOR2X1_34/B gnd NOR2X1_34/Y vdd NOR2X1
XNOR2X1_113 INVX2_102/Y NOR2X1_97/B gnd NOR2X1_113/Y vdd NOR2X1
XNOR2X1_124 INVX2_112/Y BUFX4_40/Y gnd NOR2X1_124/Y vdd NOR2X1
XNOR2X1_102 INVX2_85/Y BUFX4_41/Y gnd NOR2X1_102/Y vdd NOR2X1
XFILL_34_6_0 gnd vdd FILL
XNOR2X1_179 AOI21X1_38/Y NOR2X1_179/B gnd NOR2X1_179/Y vdd NOR2X1
XOAI21X1_608 NOR2X1_282/Y INVX2_103/Y BUFX4_122/Y gnd AOI21X1_212/C vdd OAI21X1
XNOR2X1_157 INVX2_149/Y BUFX4_217/Y gnd NOR2X1_157/Y vdd NOR2X1
XNOR2X1_168 INVX2_158/Y NOR2X1_97/B gnd NOR2X1_168/Y vdd NOR2X1
XNOR2X1_146 INVX2_132/Y NOR2X1_71/B gnd NOR2X1_146/Y vdd NOR2X1
XNOR2X1_135 INVX2_122/Y NOR2X1_76/B gnd NOR2X1_135/Y vdd NOR2X1
XOAI21X1_619 OAI21X1_619/A OAI21X1_619/B NAND2X1_272/Y gnd DFFSR_160/D vdd OAI21X1
XINVX1_15 INVX1_15/A gnd INVX1_15/Y vdd INVX1
XINVX1_26 INVX1_26/A gnd INVX1_26/Y vdd INVX1
XINVX1_37 INVX1_37/A gnd INVX1_37/Y vdd INVX1
XINVX1_48 INVX1_48/A gnd INVX1_48/Y vdd INVX1
XINVX1_59 INVX1_59/A gnd INVX1_59/Y vdd INVX1
XFILL_25_6_0 gnd vdd FILL
XFILL_0_6_0 gnd vdd FILL
XAOI21X1_260 AOI21X1_259/Y AOI21X1_260/B NOR2X1_333/Y gnd DFFSR_163/D vdd AOI21X1
XFILL_16_6_0 gnd vdd FILL
XOAI21X1_427 OAI21X1_427/A OAI21X1_427/B OAI21X1_427/C gnd DFFSR_215/D vdd OAI21X1
XOAI21X1_449 BUFX4_65/Y NAND2X1_249/Y OAI21X1_449/C gnd AOI21X1_156/B vdd OAI21X1
XOAI21X1_405 OAI21X1_405/A OAI21X1_405/B OAI21X1_401/Y gnd DFFSR_221/D vdd OAI21X1
XOAI21X1_438 BUFX4_99/Y INVX4_6/Y INVX1_123/A gnd OR2X2_14/A vdd OAI21X1
XOAI21X1_416 BUFX4_221/Y BUFX4_233/Y INVX1_40/A gnd OAI21X1_416/Y vdd OAI21X1
XDFFSR_251 OR2X2_7/B DFFSR_71/CLK DFFSR_165/R vdd DFFSR_251/D gnd vdd DFFSR
XDFFSR_240 INVX2_81/A CLKBUF1_34/A DFFSR_194/R vdd DFFSR_240/D gnd vdd DFFSR
XINVX2_80 INVX2_80/A gnd INVX2_80/Y vdd INVX2
XINVX2_91 INVX2_91/A gnd INVX2_91/Y vdd INVX2
XOAI21X1_32 BUFX4_179/Y INVX1_16/Y NAND3X1_18/Y gnd DFFSR_24/D vdd OAI21X1
XOAI21X1_54 BUFX4_181/Y INVX2_11/Y NAND3X1_29/Y gnd DFFSR_3/D vdd OAI21X1
XOAI21X1_76 NAND2X1_33/Y INVX1_21/Y DFFSR_41/Q gnd OAI21X1_76/Y vdd OAI21X1
XFILL_31_4_0 gnd vdd FILL
XOAI21X1_87 AND2X2_2/Y INVX2_20/Y NAND3X1_46/Y gnd DFFSR_37/D vdd OAI21X1
XOAI21X1_21 INVX1_11/Y BUFX4_164/Y OAI21X1_21/C gnd NAND3X1_13/B vdd OAI21X1
XOAI21X1_65 INVX1_17/Y BUFX4_5/Y OAI21X1_65/C gnd OAI21X1_65/Y vdd OAI21X1
XOAI21X1_43 INVX2_6/Y BUFX4_8/Y OAI21X1_73/C gnd OAI21X1_43/Y vdd OAI21X1
XOAI21X1_98 INVX2_25/Y BUFX4_5/Y OAI21X1_67/C gnd NAND3X1_53/B vdd OAI21X1
XOAI21X1_10 BUFX4_180/Y INVX1_5/Y NAND3X1_7/Y gnd DFFSR_29/D vdd OAI21X1
XFILL_22_4_0 gnd vdd FILL
XOAI21X1_279 AOI21X1_46/Y AND2X2_19/Y INVX8_9/Y gnd AND2X2_21/B vdd OAI21X1
XOAI21X1_268 INVX1_103/A INVX8_13/Y INVX2_48/A gnd NAND2X1_129/A vdd OAI21X1
XOAI21X1_235 NOR2X1_117/Y NOR2X1_118/Y BUFX4_184/Y gnd NAND3X1_136/C vdd OAI21X1
XOAI21X1_202 INVX8_9/A INVX1_89/A OAI21X1_202/C gnd BUFX4_45/A vdd OAI21X1
XOAI21X1_224 NOR2X1_108/Y NOR2X1_107/Y BUFX4_188/Y gnd OAI21X1_224/Y vdd OAI21X1
XOAI21X1_257 NOR2X1_158/Y NOR2X1_159/Y BUFX4_195/Y gnd OAI21X1_257/Y vdd OAI21X1
XOAI21X1_246 NOR2X1_139/Y NOR2X1_140/Y BUFX4_195/Y gnd OAI21X1_246/Y vdd OAI21X1
XOAI21X1_213 NOR2X1_85/Y NOR2X1_86/Y BUFX4_187/Y gnd NAND3X1_117/C vdd OAI21X1
XAND2X2_13 AND2X2_13/A BUFX4_187/Y gnd AND2X2_13/Y vdd AND2X2
XNAND2X1_252 INVX4_7/A AND2X2_26/A gnd AOI21X1_163/B vdd NAND2X1
XNAND2X1_241 INVX8_17/A INVX1_127/Y gnd AOI21X1_137/B vdd NAND2X1
XNAND2X1_230 INVX8_17/A AND2X2_22/A gnd NAND2X1_230/Y vdd NAND2X1
XAND2X2_24 AND2X2_24/A INVX4_8/A gnd AND2X2_24/Y vdd AND2X2
XNAND2X1_296 INVX8_22/A INVX1_150/Y gnd NAND2X1_296/Y vdd NAND2X1
XNAND2X1_285 INVX1_143/A BUFX4_62/Y gnd AOI22X1_79/C vdd NAND2X1
XFILL_5_5_0 gnd vdd FILL
XNAND2X1_263 DFFSR_172/Q BUFX4_205/Y gnd NAND2X1_263/Y vdd NAND2X1
XNAND2X1_274 INVX4_10/A INVX1_139/Y gnd AOI21X1_223/B vdd NAND2X1
XFILL_13_4_0 gnd vdd FILL
XOAI21X1_791 XNOR2X1_12/Y INVX4_5/Y OAI21X1_791/C gnd DFFSR_246/D vdd OAI21X1
XOAI21X1_780 INVX1_98/Y BUFX4_10/Y NAND2X1_328/Y gnd NAND2X1_337/B vdd OAI21X1
XDFFSR_24 INVX1_16/A CLKBUF1_37/Y DFFSR_2/R vdd DFFSR_24/D gnd vdd DFFSR
XDFFSR_35 INVX4_2/A DFFSR_5/CLK DFFSR_1/R vdd DFFSR_35/D gnd vdd DFFSR
XDFFSR_13 INVX2_5/A CLKBUF1_23/Y DFFSR_53/R vdd DFFSR_13/D gnd vdd DFFSR
XDFFSR_46 INVX8_3/A DFFSR_46/CLK DFFSR_58/R vdd DFFSR_46/D gnd vdd DFFSR
XCLKBUF1_22 CLKBUF1_54/Y gnd DFFSR_88/CLK vdd CLKBUF1
XDFFSR_68 DFFSR_68/Q DFFSR_8/CLK DFFSR_1/R vdd DFFSR_68/D gnd vdd DFFSR
XDFFSR_57 DFFSR_57/Q DFFSR_87/CLK DFFSR_58/R vdd DFFSR_57/D gnd vdd DFFSR
XCLKBUF1_11 CLKBUF1_56/Y gnd CLKBUF1_11/Y vdd CLKBUF1
XDFFSR_79 DFFSR_79/Q CLKBUF1_8/Y DFFSR_25/R vdd DFFSR_79/D gnd vdd DFFSR
XCLKBUF1_33 CLKBUF1_34/A gnd CLKBUF1_33/Y vdd CLKBUF1
XCLKBUF1_44 CLKBUF1_4/A gnd DFFSR_83/CLK vdd CLKBUF1
XCLKBUF1_55 wb_clk_i gnd CLKBUF1_55/Y vdd CLKBUF1
XCLKBUF1_66 wb_clk_i gnd CLKBUF1_34/A vdd CLKBUF1
XINVX1_107 INVX1_107/A gnd INVX1_107/Y vdd INVX1
XINVX1_118 INVX1_118/A gnd INVX1_118/Y vdd INVX1
XINVX1_129 INVX1_129/A gnd INVX1_129/Y vdd INVX1
XFILL_27_3_0 gnd vdd FILL
XFILL_2_3_0 gnd vdd FILL
XFILL_10_2_0 gnd vdd FILL
XBUFX4_246 DFFSR_44/Q gnd INVX2_18/A vdd BUFX4
XBUFX4_213 BUFX4_217/A gnd NOR2X1_97/B vdd BUFX4
XFILL_18_3_0 gnd vdd FILL
XBUFX4_202 BUFX4_200/A gnd INVX8_4/A vdd BUFX4
XBUFX4_224 INVX8_12/Y gnd BUFX4_224/Y vdd BUFX4
XNOR2X1_306 INVX1_148/Y BUFX4_63/Y gnd NOR2X1_306/Y vdd NOR2X1
XBUFX4_235 BUFX4_239/A gnd INVX8_10/A vdd BUFX4
XNOR2X1_339 BUFX4_33/Y OR2X2_20/A gnd INVX1_164/A vdd NOR2X1
XNOR2X1_328 BUFX4_229/Y NOR2X1_329/B gnd AND2X2_31/A vdd NOR2X1
XNOR2X1_317 INVX1_155/Y BUFX4_64/Y gnd NOR2X1_317/Y vdd NOR2X1
XNAND3X1_13 BUFX4_19/Y NAND3X1_13/B BUFX4_26/Y gnd OAI21X1_22/C vdd NAND3X1
XNAND3X1_46 NAND3X1_46/A BUFX4_16/Y INVX8_2/Y gnd NAND3X1_46/Y vdd NAND3X1
XNAND3X1_68 wb_adr_i[2] INVX2_39/Y INVX2_17/Y gnd OAI22X1_4/C vdd NAND3X1
XNAND3X1_35 wb_adr_i[4] INVX4_1/Y INVX2_17/Y gnd INVX8_2/A vdd NAND3X1
XNAND3X1_24 BUFX4_20/Y OAI21X1_43/Y BUFX4_27/Y gnd OAI21X1_44/C vdd NAND3X1
XNAND3X1_79 wb_adr_i[4] DFFSR_41/Q NOR2X1_3/Y gnd NAND2X1_48/B vdd NAND3X1
XNOR2X1_35 INVX2_37/A DFFSR_54/Q gnd NOR2X1_35/Y vdd NOR2X1
XNOR2X1_13 NOR2X1_13/A NOR2X1_13/B gnd NOR2X1_13/Y vdd NOR2X1
XNOR2X1_46 INVX2_29/A NOR2X1_46/B gnd NOR2X1_46/Y vdd NOR2X1
XNOR2X1_24 OR2X2_5/B DFFSR_112/Q gnd NOR2X1_24/Y vdd NOR2X1
XNAND3X1_57 AND2X2_1/B NAND3X1_57/B BUFX4_108/Y gnd NAND3X1_57/Y vdd NAND3X1
XNOR2X1_57 INVX4_3/A INVX2_48/Y gnd INVX1_88/A vdd NOR2X1
XNOR2X1_68 OR2X2_9/B OR2X2_9/A gnd NOR2X1_68/Y vdd NOR2X1
XNOR2X1_79 INVX2_64/Y BUFX4_43/Y gnd NOR2X1_79/Y vdd NOR2X1
XFILL_34_6_1 gnd vdd FILL
XNOR2X1_114 INVX2_103/Y BUFX4_45/Y gnd NOR2X1_114/Y vdd NOR2X1
XNOR2X1_147 INVX2_133/Y BUFX4_42/Y gnd NOR2X1_147/Y vdd NOR2X1
XNOR2X1_158 INVX2_150/Y NOR2X1_99/B gnd NOR2X1_158/Y vdd NOR2X1
XNOR2X1_125 INVX2_113/Y NOR2X1_87/B gnd NOR2X1_125/Y vdd NOR2X1
XNOR2X1_136 INVX2_123/Y BUFX4_40/Y gnd NOR2X1_136/Y vdd NOR2X1
XNOR2X1_103 INVX2_86/Y BUFX4_215/Y gnd NOR2X1_103/Y vdd NOR2X1
XFILL_33_1_0 gnd vdd FILL
XOAI21X1_609 INVX2_103/Y BUFX4_160/Y NAND2X1_229/Y gnd OAI21X1_609/Y vdd OAI21X1
XNOR2X1_169 INVX2_159/Y BUFX4_42/Y gnd NOR2X1_169/Y vdd NOR2X1
XFILL_16_1 gnd vdd FILL
XDFFSR_1 DFFSR_1/Q DFFSR_1/CLK DFFSR_1/R vdd DFFSR_1/D gnd vdd DFFSR
XINVX1_16 INVX1_16/A gnd INVX1_16/Y vdd INVX1
XINVX1_27 INVX1_27/A gnd INVX1_27/Y vdd INVX1
XINVX1_38 INVX1_38/A gnd INVX1_38/Y vdd INVX1
XINVX1_49 INVX1_49/A gnd INVX1_49/Y vdd INVX1
XFILL_25_6_1 gnd vdd FILL
XFILL_24_1_0 gnd vdd FILL
XNAND2X1_90 INVX2_33/A BUFX4_1/Y gnd NAND2X1_90/Y vdd NAND2X1
XFILL_0_6_1 gnd vdd FILL
XAOI21X1_261 INVX2_129/Y OR2X2_20/Y BUFX4_31/Y gnd OAI21X1_772/C vdd AOI21X1
XAOI21X1_250 NOR2X1_326/Y BUFX4_67/Y AOI21X1_250/C gnd AOI21X1_250/Y vdd AOI21X1
XFILL_7_2_0 gnd vdd FILL
XFILL_16_6_1 gnd vdd FILL
XFILL_15_1_0 gnd vdd FILL
XDFFSR_252 XOR2X1_3/A CLKBUF1_27/Y DFFSR_165/R vdd DFFSR_252/D gnd vdd DFFSR
XOAI21X1_428 BUFX4_66/Y OR2X2_12/Y AOI21X1_141/Y gnd OAI21X1_428/Y vdd OAI21X1
XDFFSR_230 INVX2_77/A CLKBUF1_1/Y DFFSR_203/R vdd DFFSR_230/D gnd vdd DFFSR
XOAI21X1_417 NOR2X1_226/Y INVX2_158/Y BUFX4_51/Y gnd AOI21X1_136/C vdd OAI21X1
XDFFSR_241 INVX2_150/A DFFSR_46/CLK DFFSR_236/R vdd DFFSR_241/D gnd vdd DFFSR
XOAI21X1_439 BUFX4_65/Y OR2X2_14/Y OAI21X1_439/C gnd AOI21X1_153/B vdd OAI21X1
XOAI21X1_406 BUFX4_221/Y BUFX4_233/Y INVX1_46/A gnd OAI21X1_410/C vdd OAI21X1
XINVX2_92 INVX1_35/A gnd INVX2_92/Y vdd INVX2
XINVX2_81 INVX2_81/A gnd INVX2_81/Y vdd INVX2
XINVX2_70 INVX1_50/A gnd INVX2_70/Y vdd INVX2
XOAI21X1_11 INVX1_6/Y BUFX4_72/Y NAND2X1_6/Y gnd NAND3X1_8/B vdd OAI21X1
XOAI21X1_77 AND2X2_2/Y OAI21X1_76/Y NAND3X1_41/Y gnd DFFSR_41/D vdd OAI21X1
XFILL_31_4_1 gnd vdd FILL
XOAI21X1_22 BUFX4_179/Y INVX1_11/Y OAI21X1_22/C gnd DFFSR_19/D vdd OAI21X1
XOAI21X1_88 INVX2_21/Y BUFX4_84/Y OAI21X1_59/C gnd NAND3X1_47/A vdd OAI21X1
XOAI21X1_55 INVX2_12/Y BUFX4_86/Y NAND2X1_28/Y gnd NAND3X1_30/B vdd OAI21X1
XOAI21X1_66 AND2X2_2/Y INVX1_17/Y NAND3X1_36/Y gnd DFFSR_42/D vdd OAI21X1
XOAI21X1_33 INVX2_1/Y BUFX4_6/Y OAI21X1_33/C gnd OAI21X1_33/Y vdd OAI21X1
XOAI21X1_44 BUFX4_182/Y INVX2_6/Y OAI21X1_44/C gnd DFFSR_14/D vdd OAI21X1
XOAI21X1_99 AND2X2_3/Y INVX2_25/Y OAI21X1_99/C gnd DFFSR_57/D vdd OAI21X1
XOAI21X1_203 BUFX4_245/Y INVX1_89/Y OAI21X1_203/C gnd BUFX4_217/A vdd OAI21X1
XFILL_22_4_1 gnd vdd FILL
XOAI21X1_258 NOR2X1_160/Y NOR2X1_161/Y AND2X2_15/B gnd NAND3X1_160/C vdd OAI21X1
XOAI21X1_269 AND2X2_9/Y NOR2X1_47/Y BUFX4_112/Y gnd AOI21X1_33/B vdd OAI21X1
XAND2X2_25 AND2X2_25/A INVX4_8/A gnd AND2X2_25/Y vdd AND2X2
XOAI21X1_225 NOR2X1_110/Y NOR2X1_109/Y BUFX4_194/Y gnd NAND3X1_130/B vdd OAI21X1
XOAI21X1_236 NOR2X1_119/Y NOR2X1_120/Y BUFX4_195/Y gnd OAI21X1_236/Y vdd OAI21X1
XOAI21X1_247 AND2X2_17/Y NOR2X1_141/Y BUFX4_187/Y gnd OAI21X1_247/Y vdd OAI21X1
XOAI21X1_214 NOR2X1_87/Y NOR2X1_88/Y AND2X2_16/B gnd OAI21X1_214/Y vdd OAI21X1
XAND2X2_14 AND2X2_14/A AND2X2_16/B gnd AND2X2_14/Y vdd AND2X2
XNAND2X1_264 INVX2_54/A BUFX4_204/Y gnd NAND2X1_264/Y vdd NAND2X1
XNAND2X1_242 BUFX4_83/Y wb_dat_i[4] gnd NAND2X1_242/Y vdd NAND2X1
XNAND2X1_253 INVX4_7/A AND2X2_27/A gnd AOI21X1_170/B vdd NAND2X1
XNAND2X1_220 INVX1_111/A NOR2X1_189/Y gnd INVX1_128/A vdd NAND2X1
XNAND2X1_286 INVX1_144/A BUFX4_62/Y gnd AOI22X1_80/C vdd NAND2X1
XFILL_5_5_1 gnd vdd FILL
XNAND2X1_231 wb_dat_i[14] BUFX4_11/Y gnd NAND2X1_231/Y vdd NAND2X1
XNAND2X1_275 INVX1_49/A BUFX4_203/Y gnd NAND2X1_275/Y vdd NAND2X1
XFILL_29_0_0 gnd vdd FILL
XNAND2X1_297 BUFX4_208/Y NAND2X1_297/B gnd OAI21X1_683/C vdd NAND2X1
XFILL_4_0_0 gnd vdd FILL
XFILL_13_4_1 gnd vdd FILL
XOAI21X1_792 OR2X2_8/B INVX4_11/A BUFX4_101/Y gnd OAI22X1_42/D vdd OAI21X1
XOAI21X1_781 INVX1_163/A INVX1_98/A BUFX4_117/Y gnd OAI21X1_781/Y vdd OAI21X1
XOAI21X1_770 INVX2_123/Y BUFX4_9/Y NAND2X1_328/Y gnd AOI21X1_259/B vdd OAI21X1
XDFFSR_36 INVX4_3/A DFFSR_36/CLK DFFSR_1/R vdd DFFSR_36/D gnd vdd DFFSR
XDFFSR_69 BUFX2_40/A DFFSR_9/CLK DFFSR_9/R vdd DFFSR_69/D gnd vdd DFFSR
XDFFSR_47 OR2X2_2/B DFFSR_47/CLK DFFSR_53/R vdd DFFSR_47/D gnd vdd DFFSR
XDFFSR_14 INVX2_6/A CLKBUF1_55/Y DFFSR_53/R vdd DFFSR_14/D gnd vdd DFFSR
XDFFSR_25 INVX1_1/A CLKBUF1_34/Y DFFSR_25/R vdd DFFSR_25/D gnd vdd DFFSR
XDFFSR_58 INVX2_26/A DFFSR_28/CLK DFFSR_58/R vdd DFFSR_58/D gnd vdd DFFSR
XCLKBUF1_12 CLKBUF1_12/A gnd CLKBUF1_12/Y vdd CLKBUF1
XCLKBUF1_23 CLKBUF1_55/Y gnd CLKBUF1_23/Y vdd CLKBUF1
XCLKBUF1_56 wb_clk_i gnd CLKBUF1_56/Y vdd CLKBUF1
XCLKBUF1_34 CLKBUF1_34/A gnd CLKBUF1_34/Y vdd CLKBUF1
XCLKBUF1_45 CLKBUF1_34/A gnd CLKBUF1_45/Y vdd CLKBUF1
XCLKBUF1_67 wb_clk_i gnd CLKBUF1_5/A vdd CLKBUF1
XINVX1_108 INVX1_108/A gnd INVX1_108/Y vdd INVX1
XINVX1_119 BUFX2_2/A gnd INVX1_119/Y vdd INVX1
XFILL_4_1 gnd vdd FILL
XFILL_27_3_1 gnd vdd FILL
XFILL_2_3_1 gnd vdd FILL
XFILL_10_2_1 gnd vdd FILL
XBUFX4_247 DFFSR_44/Q gnd INVX8_9/A vdd BUFX4
XNOR2X1_307 BUFX4_32/Y OR2X2_17/A gnd INVX1_149/A vdd NOR2X1
XBUFX4_225 BUFX4_228/A gnd OAI22X1_9/A vdd BUFX4
XFILL_18_3_1 gnd vdd FILL
XBUFX4_203 BUFX4_211/A gnd BUFX4_203/Y vdd BUFX4
XBUFX4_214 BUFX4_217/A gnd NOR2X1_99/B vdd BUFX4
XNOR2X1_318 OR2X2_18/B NOR2X1_300/B gnd INVX1_156/A vdd NOR2X1
XNOR2X1_329 INVX4_8/Y NOR2X1_329/B gnd NOR2X1_329/Y vdd NOR2X1
XBUFX4_236 BUFX4_239/A gnd MUX2X1_1/S vdd BUFX4
XNAND3X1_14 BUFX4_19/Y NAND3X1_14/B BUFX4_26/Y gnd NAND3X1_14/Y vdd NAND3X1
XNOR2X1_58 NOR2X1_56/Y INVX1_88/A gnd NOR2X1_58/Y vdd NOR2X1
XNOR2X1_47 OR2X2_8/A OR2X2_8/B gnd NOR2X1_47/Y vdd NOR2X1
XNAND3X1_69 wb_adr_i[3] DFFSR_180/Q NOR2X1_4/Y gnd NAND3X1_69/Y vdd NAND3X1
XNAND3X1_47 NAND3X1_47/A BUFX4_19/Y INVX8_2/Y gnd NAND3X1_47/Y vdd NAND3X1
XNOR2X1_69 INVX2_55/Y NOR2X1_97/B gnd NOR2X1_69/Y vdd NOR2X1
XNAND3X1_36 OAI21X1_65/Y BUFX4_18/Y INVX8_2/Y gnd NAND3X1_36/Y vdd NAND3X1
XNAND3X1_25 BUFX4_18/Y OAI21X1_45/Y BUFX4_27/Y gnd NAND3X1_25/Y vdd NAND3X1
XNOR2X1_36 DFFSR_51/Q INVX2_36/A gnd NOR2X1_36/Y vdd NOR2X1
XNOR2X1_25 OR2X2_6/B DFFSR_114/Q gnd INVX1_78/A vdd NOR2X1
XNOR2X1_14 NOR2X1_14/A NOR2X1_14/B gnd NOR2X1_14/Y vdd NOR2X1
XNAND3X1_58 AND2X2_1/B NAND3X1_58/B BUFX4_108/Y gnd NAND3X1_58/Y vdd NAND3X1
XFILL_33_1_1 gnd vdd FILL
XNOR2X1_115 INVX2_104/Y NOR2X1_97/B gnd NOR2X1_115/Y vdd NOR2X1
XNOR2X1_148 INVX2_134/Y NOR2X1_71/B gnd NOR2X1_148/Y vdd NOR2X1
XNOR2X1_159 INVX2_151/Y BUFX4_43/Y gnd NOR2X1_159/Y vdd NOR2X1
XNOR2X1_137 INVX2_124/Y NOR2X1_87/B gnd NOR2X1_137/Y vdd NOR2X1
XNOR2X1_126 INVX1_97/Y BUFX4_40/Y gnd NOR2X1_126/Y vdd NOR2X1
XMUX2X1_10 wb_dat_i[10] INVX1_94/A BUFX4_11/Y gnd MUX2X1_10/Y vdd MUX2X1
XNOR2X1_104 INVX2_87/Y BUFX4_41/Y gnd NOR2X1_104/Y vdd NOR2X1
XDFFSR_2 DFFSR_2/Q DFFSR_2/CLK DFFSR_2/R vdd DFFSR_2/D gnd vdd DFFSR
XFILL_16_2 gnd vdd FILL
XINVX1_39 INVX1_39/A gnd INVX1_39/Y vdd INVX1
XINVX1_28 INVX1_28/A gnd INVX1_28/Y vdd INVX1
XINVX1_17 INVX1_17/A gnd INVX1_17/Y vdd INVX1
XNAND2X1_80 AND2X2_4/A AND2X2_4/B gnd NOR3X1_2/A vdd NAND2X1
XNAND2X1_91 OR2X2_2/A BUFX4_1/Y gnd NAND2X1_91/Y vdd NAND2X1
XFILL_24_1_1 gnd vdd FILL
XAOI21X1_240 NOR2X1_293/Y BUFX4_58/Y OAI21X1_640/Y gnd OAI21X1_643/A vdd AOI21X1
XAOI21X1_262 BUFX4_31/Y AOI21X1_262/B BUFX4_203/Y gnd AOI21X1_262/Y vdd AOI21X1
XAOI21X1_251 NOR2X1_327/Y BUFX4_59/Y AOI21X1_251/C gnd OAI21X1_750/A vdd AOI21X1
XFILL_7_2_1 gnd vdd FILL
XFILL_15_1_1 gnd vdd FILL
XNAND3X1_200 DFFSR_133/Q OAI21X1_287/Y NAND3X1_198/Y gnd OAI21X1_295/C vdd NAND3X1
XDFFSR_253 NOR2X1_50/A DFFSR_88/CLK DFFSR_165/R vdd DFFSR_253/D gnd vdd DFFSR
XOAI21X1_429 INVX2_75/Y BUFX4_80/Y NAND2X1_244/Y gnd OAI21X1_429/Y vdd OAI21X1
XOAI21X1_418 INVX2_158/Y BUFX4_82/Y NAND2X1_240/Y gnd OAI21X1_419/B vdd OAI21X1
XDFFSR_231 AOI22X1_8/C CLKBUF1_50/Y DFFSR_203/R vdd DFFSR_231/D gnd vdd DFFSR
XDFFSR_242 INVX2_65/A DFFSR_92/CLK DFFSR_236/R vdd DFFSR_242/D gnd vdd DFFSR
XDFFSR_220 INVX1_46/A CLKBUF1_33/Y DFFSR_203/R vdd DFFSR_220/D gnd vdd DFFSR
XOAI21X1_407 NOR2X1_224/Y INVX2_99/Y BUFX4_54/Y gnd AOI21X1_134/C vdd OAI21X1
XINVX2_60 INVX2_60/A gnd INVX2_60/Y vdd INVX2
XINVX2_93 INVX1_37/A gnd INVX2_93/Y vdd INVX2
XINVX2_82 INVX2_82/A gnd INVX2_82/Y vdd INVX2
XINVX2_71 INVX1_51/A gnd INVX2_71/Y vdd INVX2
XOAI21X1_23 INVX1_12/Y NAND2X1_9/B NAND2X1_12/Y gnd NAND3X1_14/B vdd OAI21X1
XOAI21X1_34 BUFX4_183/Y INVX2_1/Y OAI21X1_34/C gnd DFFSR_9/D vdd OAI21X1
XOAI21X1_45 INVX2_7/Y BUFX4_10/Y OAI21X1_45/C gnd OAI21X1_45/Y vdd OAI21X1
XOAI21X1_12 BUFX4_180/Y INVX1_6/Y NAND3X1_8/Y gnd DFFSR_30/D vdd OAI21X1
XOAI21X1_89 AND2X2_2/Y INVX2_21/Y NAND3X1_47/Y gnd DFFSR_38/D vdd OAI21X1
XOAI21X1_78 INVX1_22/Y BUFX4_79/Y NAND2X1_25/Y gnd NAND3X1_42/A vdd OAI21X1
XOAI21X1_56 BUFX4_183/Y INVX2_12/Y OAI21X1_56/C gnd DFFSR_4/D vdd OAI21X1
XOAI21X1_67 INVX1_18/Y BUFX4_6/Y OAI21X1_67/C gnd OAI21X1_67/Y vdd OAI21X1
XOAI21X1_226 NOR2X1_112/Y NOR2X1_111/Y BUFX4_185/Y gnd NAND3X1_130/C vdd OAI21X1
XOAI21X1_204 XNOR2X1_6/Y INVX8_9/Y OAI21X1_204/C gnd BUFX4_185/A vdd OAI21X1
XOAI21X1_237 NOR2X1_121/Y NOR2X1_122/Y AND2X2_15/B gnd OAI21X1_237/Y vdd OAI21X1
XOAI21X1_215 NOR2X1_89/Y NOR2X1_90/Y BUFX4_187/Y gnd NAND3X1_118/C vdd OAI21X1
XAND2X2_26 AND2X2_26/A INVX4_8/A gnd AND2X2_26/Y vdd AND2X2
XOAI21X1_248 NOR2X1_142/Y NOR2X1_143/Y BUFX4_197/Y gnd OAI21X1_248/Y vdd OAI21X1
XAND2X2_15 AND2X2_15/A AND2X2_15/B gnd AND2X2_15/Y vdd AND2X2
XOAI21X1_259 NOR2X1_162/Y NOR2X1_163/Y BUFX4_197/Y gnd NAND3X1_161/B vdd OAI21X1
XFILL_29_0_1 gnd vdd FILL
XNAND2X1_243 BUFX4_85/Y wb_dat_i[3] gnd NAND2X1_243/Y vdd NAND2X1
XNAND2X1_221 INVX8_14/A INVX1_128/Y gnd NAND2X1_221/Y vdd NAND2X1
XNAND2X1_265 INVX4_9/A NOR2X1_276/Y gnd NAND2X1_265/Y vdd NAND2X1
XNAND2X1_298 INVX8_22/A INVX1_151/Y gnd OAI21X1_682/B vdd NAND2X1
XNAND2X1_232 BUFX4_5/Y wb_dat_i[13] gnd NAND2X1_232/Y vdd NAND2X1
XFILL_4_0_1 gnd vdd FILL
XNAND2X1_210 MUX2X1_7/S wb_dat_i[25] gnd OAI21X1_458/C vdd NAND2X1
XNAND2X1_287 INVX1_145/A BUFX4_62/Y gnd AOI22X1_81/C vdd NAND2X1
XNAND2X1_254 INVX4_8/A INVX1_131/Y gnd AOI21X1_172/B vdd NAND2X1
XNAND2X1_276 INVX4_10/A INVX1_140/Y gnd OAI21X1_628/B vdd NAND2X1
XOAI21X1_793 NAND2X1_104/Y INVX4_11/Y BUFX4_101/Y gnd OAI22X1_43/C vdd OAI21X1
XOAI21X1_771 BUFX4_98/Y INVX8_11/Y AND2X2_32/A gnd OR2X2_20/A vdd OAI21X1
XOAI21X1_760 BUFX4_59/Y NAND2X1_332/Y OAI21X1_760/C gnd AOI21X1_255/B vdd OAI21X1
XOAI21X1_782 NOR2X1_338/Y OAI21X1_781/Y OAI21X1_782/C gnd DFFSR_131/D vdd OAI21X1
XDFFSR_37 INVX2_49/A DFFSR_82/CLK DFFSR_2/R vdd DFFSR_37/D gnd vdd DFFSR
XDFFSR_48 INVX2_32/A DFFSR_3/CLK DFFSR_9/R vdd DFFSR_48/D gnd vdd DFFSR
XDFFSR_15 INVX2_7/A CLKBUF1_7/A DFFSR_9/R vdd DFFSR_15/D gnd vdd DFFSR
XDFFSR_59 INVX2_27/A DFFSR_59/CLK DFFSR_58/R vdd DFFSR_59/D gnd vdd DFFSR
XDFFSR_26 INVX1_2/A DFFSR_26/CLK DFFSR_25/R vdd DFFSR_26/D gnd vdd DFFSR
XCLKBUF1_46 CLKBUF1_46/A gnd DFFSR_82/CLK vdd CLKBUF1
XCLKBUF1_35 CLKBUF1_7/A gnd CLKBUF1_35/Y vdd CLKBUF1
XCLKBUF1_13 CLKBUF1_5/A gnd CLKBUF1_13/Y vdd CLKBUF1
XCLKBUF1_57 wb_clk_i gnd CLKBUF1_38/A vdd CLKBUF1
XCLKBUF1_24 CLKBUF1_34/A gnd CLKBUF1_24/Y vdd CLKBUF1
XINVX1_109 XOR2X1_4/Y gnd INVX1_109/Y vdd INVX1
XOAI21X1_590 BUFX4_98/Y INVX8_11/Y AND2X2_26/A gnd OR2X2_16/A vdd OAI21X1
XFILL_4_2 gnd vdd FILL
XNOR2X1_308 BUFX4_28/Y OR2X2_16/A gnd NOR2X1_308/Y vdd NOR2X1
XBUFX4_248 DFFSR_44/Q gnd BUFX4_248/Y vdd BUFX4
XBUFX4_204 BUFX4_211/A gnd BUFX4_204/Y vdd BUFX4
XBUFX4_237 BUFX4_239/A gnd BUFX4_237/Y vdd BUFX4
XBUFX4_215 BUFX4_217/A gnd BUFX4_215/Y vdd BUFX4
XBUFX4_226 BUFX4_228/A gnd BUFX4_226/Y vdd BUFX4
XNOR2X1_319 OR2X2_18/B NOR2X1_301/B gnd INVX1_157/A vdd NOR2X1
XFILL_20_5_0 gnd vdd FILL
XNAND3X1_15 BUFX4_19/Y NAND3X1_15/B BUFX4_26/Y gnd OAI21X1_26/C vdd NAND3X1
XNAND3X1_48 OAI21X1_90/Y BUFX4_16/Y INVX8_2/Y gnd NAND3X1_48/Y vdd NAND3X1
XNAND3X1_37 OAI21X1_67/Y BUFX4_18/Y INVX8_2/Y gnd OAI21X1_68/C vdd NAND3X1
XNAND3X1_26 AND2X2_1/B NAND3X1_26/B BUFX4_23/Y gnd OAI21X1_48/C vdd NAND3X1
XNOR2X1_48 INVX2_48/A NOR2X1_48/B gnd INVX1_86/A vdd NOR2X1
XNOR2X1_59 NOR2X1_58/Y AND2X2_10/A gnd NOR2X1_59/Y vdd NOR2X1
XFILL_28_6_0 gnd vdd FILL
XNAND3X1_59 AND2X2_2/B NAND3X1_59/B BUFX4_106/Y gnd NAND3X1_59/Y vdd NAND3X1
XNOR2X1_15 NOR2X1_15/A NOR2X1_15/B gnd NOR2X1_15/Y vdd NOR2X1
XNOR2X1_37 INVX2_33/A INVX2_32/A gnd NOR2X1_37/Y vdd NOR2X1
XFILL_3_6_0 gnd vdd FILL
XNOR2X1_26 NOR3X1_2/B INVX1_77/A gnd NOR2X1_26/Y vdd NOR2X1
XFILL_11_5_0 gnd vdd FILL
XFILL_19_6_0 gnd vdd FILL
XMUX2X1_11 wb_dat_i[31] AND2X2_17/B MUX2X1_6/S gnd MUX2X1_11/Y vdd MUX2X1
XNOR2X1_116 INVX2_105/Y BUFX4_44/Y gnd NOR2X1_116/Y vdd NOR2X1
XNOR2X1_149 INVX2_135/Y BUFX4_42/Y gnd NOR2X1_149/Y vdd NOR2X1
XNOR2X1_127 INVX2_114/Y BUFX4_215/Y gnd NOR2X1_127/Y vdd NOR2X1
XNOR2X1_105 INVX2_88/Y BUFX4_46/Y gnd NOR2X1_105/Y vdd NOR2X1
XNOR2X1_138 INVX1_98/Y BUFX4_40/Y gnd NOR2X1_138/Y vdd NOR2X1
XDFFSR_3 DFFSR_3/Q DFFSR_3/CLK DFFSR_2/R vdd DFFSR_3/D gnd vdd DFFSR
XFILL_16_3 gnd vdd FILL
XINVX1_29 INVX1_29/A gnd INVX1_29/Y vdd INVX1
XINVX1_18 DFFSR_43/Q gnd INVX1_18/Y vdd INVX1
XNAND2X1_70 INVX1_93/A BUFX4_192/Y gnd NAND3X1_96/B vdd NAND2X1
XNAND2X1_81 NOR2X1_27/Y NOR2X1_31/Y gnd OAI22X1_41/A vdd NAND2X1
XNAND2X1_92 INVX2_36/A BUFX4_1/Y gnd NAND2X1_92/Y vdd NAND2X1
XAOI21X1_241 NOR2X1_294/Y BUFX4_61/Y AOI21X1_241/C gnd AOI21X1_241/Y vdd AOI21X1
XAOI21X1_230 INVX2_58/Y OR2X2_17/Y BUFX4_33/Y gnd AOI21X1_230/Y vdd AOI21X1
XAOI21X1_252 AND2X2_31/Y BUFX4_63/Y AOI21X1_252/C gnd OAI21X1_754/A vdd AOI21X1
XAOI21X1_263 AOI21X1_262/Y OAI21X1_772/Y NOR2X1_334/Y gnd DFFSR_171/D vdd AOI21X1
XNAND3X1_201 DFFSR_121/Q OAI21X1_287/Y NAND3X1_198/Y gnd OAI21X1_296/C vdd NAND3X1
XFILL_34_4_0 gnd vdd FILL
XOAI21X1_408 INVX2_99/Y BUFX4_8/Y NAND2X1_238/Y gnd OAI21X1_408/Y vdd OAI21X1
XOAI21X1_419 BUFX4_51/Y OAI21X1_419/B BUFX4_243/Y gnd OAI21X1_420/B vdd OAI21X1
XDFFSR_232 INVX2_89/A CLKBUF1_48/Y BUFX4_130/Y vdd DFFSR_232/D gnd vdd DFFSR
XDFFSR_243 DFFSR_243/Q CLKBUF1_11/Y DFFSR_236/R vdd DFFSR_243/D gnd vdd DFFSR
XDFFSR_210 INVX2_66/A CLKBUF1_56/Y DFFSR_236/R vdd DFFSR_210/D gnd vdd DFFSR
XDFFSR_221 INVX1_48/A CLKBUF1_32/Y DFFSR_203/R vdd DFFSR_221/D gnd vdd DFFSR
XFILL_25_4_0 gnd vdd FILL
XFILL_0_4_0 gnd vdd FILL
XFILL_8_5_0 gnd vdd FILL
XINVX2_50 INVX2_50/A gnd INVX2_50/Y vdd INVX2
XINVX2_94 INVX2_94/A gnd INVX2_94/Y vdd INVX2
XINVX2_83 INVX2_83/A gnd INVX2_83/Y vdd INVX2
XINVX2_72 INVX2_72/A gnd INVX2_72/Y vdd INVX2
XINVX2_61 INVX2_61/A gnd INVX2_61/Y vdd INVX2
XOAI21X1_24 BUFX4_179/Y INVX1_12/Y NAND3X1_14/Y gnd DFFSR_20/D vdd OAI21X1
XOAI21X1_57 INVX2_13/Y BUFX4_80/Y OAI21X1_86/C gnd NAND3X1_31/B vdd OAI21X1
XOAI21X1_46 BUFX4_183/Y INVX2_7/Y NAND3X1_25/Y gnd DFFSR_15/D vdd OAI21X1
XOAI21X1_68 AND2X2_2/Y INVX1_18/Y OAI21X1_68/C gnd DFFSR_43/D vdd OAI21X1
XOAI21X1_35 INVX2_2/Y BUFX4_8/Y OAI21X1_65/C gnd NAND3X1_20/B vdd OAI21X1
XFILL_16_4_0 gnd vdd FILL
XOAI21X1_13 INVX1_7/Y MUX2X1_6/S NAND2X1_7/Y gnd NAND3X1_9/B vdd OAI21X1
XOAI21X1_79 AND2X2_2/Y INVX1_22/Y OAI21X1_79/C gnd DFFSR_33/D vdd OAI21X1
XOAI21X1_216 NOR2X1_91/Y NOR2X1_92/Y BUFX4_184/Y gnd NAND3X1_120/B vdd OAI21X1
XOAI21X1_205 NOR2X1_69/Y NOR2X1_70/Y BUFX4_185/Y gnd NAND3X1_110/C vdd OAI21X1
XOAI21X1_249 NOR2X1_144/Y NOR2X1_145/Y BUFX4_185/Y gnd NAND3X1_151/C vdd OAI21X1
XOAI21X1_227 INVX1_120/A INVX8_10/A OAI21X1_227/C gnd AND2X2_13/A vdd OAI21X1
XOAI21X1_238 NOR2X1_123/Y NOR2X1_124/Y BUFX4_195/Y gnd OAI21X1_238/Y vdd OAI21X1
XAND2X2_27 AND2X2_27/A INVX4_8/A gnd AND2X2_27/Y vdd AND2X2
XNAND2X1_200 AOI22X1_75/Y AOI22X1_76/Y gnd NAND2X1_200/Y vdd NAND2X1
XAND2X2_16 AND2X2_16/A AND2X2_16/B gnd AND2X2_16/Y vdd AND2X2
XNAND2X1_211 INVX1_126/Y NOR2X1_191/Y gnd NOR2X1_224/A vdd NAND2X1
XNAND2X1_222 BUFX4_160/Y wb_dat_i[19] gnd NAND2X1_222/Y vdd NAND2X1
XNAND2X1_277 INVX1_38/A BUFX4_211/Y gnd NAND2X1_277/Y vdd NAND2X1
XNAND2X1_244 BUFX4_79/Y wb_dat_i[2] gnd NAND2X1_244/Y vdd NAND2X1
XNAND2X1_299 INVX8_22/A NOR2X1_309/Y gnd NAND2X1_299/Y vdd NAND2X1
XNAND2X1_266 INVX4_9/A NOR2X1_278/Y gnd NAND2X1_266/Y vdd NAND2X1
XNAND2X1_233 BUFX4_7/Y wb_dat_i[12] gnd OAI21X1_699/C vdd NAND2X1
XNAND2X1_288 BUFX4_205/Y OAI21X1_660/Y gnd OAI21X1_662/C vdd NAND2X1
XNAND2X1_255 INVX4_8/A INVX1_133/Y gnd AOI21X1_176/B vdd NAND2X1
XOAI21X1_794 INVX1_107/A INVX4_11/Y BUFX4_101/Y gnd OAI22X1_44/C vdd OAI21X1
XOAI21X1_783 INVX1_164/Y INVX8_22/Y INVX2_131/Y gnd OAI21X1_784/C vdd OAI21X1
XOAI21X1_761 INVX2_130/Y BUFX4_163/Y NAND2X1_330/Y gnd OAI21X1_762/B vdd OAI21X1
XOAI21X1_772 BUFX4_64/Y OR2X2_20/Y OAI21X1_772/C gnd OAI21X1_772/Y vdd OAI21X1
XOAI21X1_750 OAI21X1_750/A OAI21X1_750/B OAI21X1_746/Y gnd DFFSR_235/D vdd OAI21X1
XFILL_31_2_0 gnd vdd FILL
XDFFSR_38 INVX2_50/A DFFSR_83/CLK DFFSR_1/R vdd DFFSR_38/D gnd vdd DFFSR
XDFFSR_49 INVX2_33/A CLKBUF1_7/Y DFFSR_7/R vdd DFFSR_49/D gnd vdd DFFSR
XDFFSR_27 INVX1_3/A CLKBUF1_28/Y DFFSR_25/R vdd DFFSR_27/D gnd vdd DFFSR
XDFFSR_16 INVX2_8/A DFFSR_46/CLK DFFSR_95/R vdd DFFSR_16/D gnd vdd DFFSR
XCLKBUF1_36 CLKBUF1_46/A gnd DFFSR_85/CLK vdd CLKBUF1
XCLKBUF1_47 CLKBUF1_5/A gnd DFFSR_7/CLK vdd CLKBUF1
XCLKBUF1_58 wb_clk_i gnd CLKBUF1_32/A vdd CLKBUF1
XCLKBUF1_14 CLKBUF1_5/A gnd DFFSR_47/CLK vdd CLKBUF1
XCLKBUF1_25 DFFSR_59/CLK gnd DFFSR_87/CLK vdd CLKBUF1
XFILL_22_2_0 gnd vdd FILL
XBUFX4_90 INVX8_8/Y gnd BUFX4_90/Y vdd BUFX4
XFILL_5_3_0 gnd vdd FILL
XFILL_13_2_0 gnd vdd FILL
XOAI21X1_591 BUFX4_58/Y OR2X2_16/Y OAI21X1_591/C gnd AOI21X1_203/B vdd OAI21X1
XOAI21X1_580 BUFX4_99/Y INVX8_11/Y INVX1_134/A gnd INVX1_140/A vdd OAI21X1
XBUFX4_227 BUFX4_228/A gnd INVX8_6/A vdd BUFX4
XBUFX4_216 BUFX4_217/A gnd NOR2X1_76/B vdd BUFX4
XBUFX4_205 BUFX4_211/A gnd BUFX4_205/Y vdd BUFX4
XNOR2X1_309 BUFX4_32/Y NOR2X1_280/B gnd NOR2X1_309/Y vdd NOR2X1
XBUFX4_238 BUFX4_239/A gnd BUFX4_238/Y vdd BUFX4
XFILL_20_5_1 gnd vdd FILL
XNAND3X1_16 BUFX4_19/Y NAND3X1_16/B BUFX4_26/Y gnd OAI21X1_28/C vdd NAND3X1
XNAND3X1_27 BUFX4_16/Y OAI21X1_49/Y BUFX4_24/Y gnd OAI21X1_50/C vdd NAND3X1
XNAND3X1_49 OAI21X1_92/Y BUFX4_15/Y INVX8_2/Y gnd OAI21X1_93/C vdd NAND3X1
XNAND3X1_38 OAI21X1_69/Y BUFX4_18/Y INVX8_2/Y gnd NAND3X1_38/Y vdd NAND3X1
XNOR2X1_49 XOR2X1_3/A OR2X2_7/Y gnd INVX1_79/A vdd NOR2X1
XFILL_28_6_1 gnd vdd FILL
XFILL_27_1_0 gnd vdd FILL
XNOR2X1_38 OR2X2_2/Y NOR2X1_38/B gnd NOR2X1_38/Y vdd NOR2X1
XNOR2X1_16 NOR2X1_16/A NOR2X1_16/B gnd NOR2X1_16/Y vdd NOR2X1
XFILL_3_6_1 gnd vdd FILL
XFILL_2_1_0 gnd vdd FILL
XNOR2X1_27 OR2X2_4/A OR2X2_4/B gnd NOR2X1_27/Y vdd NOR2X1
XFILL_10_0_0 gnd vdd FILL
XFILL_11_5_1 gnd vdd FILL
XFILL_19_6_1 gnd vdd FILL
XFILL_18_1_0 gnd vdd FILL
XNOR2X1_106 INVX2_89/Y BUFX4_215/Y gnd NOR2X1_106/Y vdd NOR2X1
XNOR2X1_117 INVX2_106/Y BUFX4_217/Y gnd NOR2X1_117/Y vdd NOR2X1
XNOR2X1_128 INVX2_115/Y BUFX4_46/Y gnd NOR2X1_128/Y vdd NOR2X1
XNOR2X1_139 INVX2_125/Y NOR2X1_99/B gnd NOR2X1_139/Y vdd NOR2X1
XDFFSR_4 DFFSR_4/Q CLKBUF1_7/Y DFFSR_1/R vdd DFFSR_4/D gnd vdd DFFSR
XINVX1_19 INVX1_19/A gnd INVX1_19/Y vdd INVX1
XNAND2X1_60 DFFSR_132/Q AOI21X1_1/B gnd NAND3X1_86/A vdd NAND2X1
XNAND2X1_82 NOR2X1_34/Y NOR2X1_38/Y gnd NAND2X1_82/Y vdd NAND2X1
XNAND2X1_93 AND2X2_4/B NOR2X1_41/Y gnd AND2X2_7/B vdd NAND2X1
XNAND2X1_71 INVX1_96/A BUFX4_192/Y gnd NAND3X1_97/A vdd NAND2X1
XAOI21X1_242 NOR2X1_295/Y BUFX4_61/Y AOI21X1_242/C gnd OAI21X1_651/A vdd AOI21X1
XAOI21X1_231 BUFX4_33/Y AOI21X1_231/B INVX8_21/A gnd AOI21X1_231/Y vdd AOI21X1
XAOI21X1_264 NOR2X1_335/Y BUFX4_60/Y AOI21X1_264/C gnd OAI21X1_777/A vdd AOI21X1
XAOI21X1_253 NOR2X1_329/Y BUFX4_57/Y AOI21X1_253/C gnd OAI21X1_759/A vdd AOI21X1
XAOI21X1_220 INVX2_112/Y AOI21X1_220/B BUFX4_30/Y gnd OAI21X1_620/C vdd AOI21X1
XAOI22X1_80 BUFX4_212/Y MUX2X1_7/Y AOI22X1_80/C AOI22X1_80/D gnd DFFSR_143/D vdd AOI22X1
XNAND3X1_202 NAND3X1_202/A OAI21X1_300/Y AOI22X1_49/Y gnd AOI22X1_50/C vdd NAND3X1
XFILL_34_4_1 gnd vdd FILL
XDFFSR_200 INVX2_91/A CLKBUF1_1/Y DFFSR_203/R vdd DFFSR_200/D gnd vdd DFFSR
XOAI21X1_409 BUFX4_54/Y OAI21X1_408/Y BUFX4_243/Y gnd OAI21X1_410/B vdd OAI21X1
XDFFSR_244 BUFX2_1/A CLKBUF1_5/Y DFFSR_137/R vdd DFFSR_244/D gnd vdd DFFSR
XDFFSR_233 DFFSR_233/Q CLKBUF1_42/Y DFFSR_203/R vdd DFFSR_233/D gnd vdd DFFSR
XDFFSR_222 INVX1_50/A CLKBUF1_26/Y DFFSR_236/R vdd DFFSR_222/D gnd vdd DFFSR
XDFFSR_211 INVX2_127/A DFFSR_46/CLK DFFSR_194/R vdd DFFSR_211/D gnd vdd DFFSR
XFILL_25_4_1 gnd vdd FILL
XFILL_0_4_1 gnd vdd FILL
XINVX2_51 OR2X2_7/B gnd INVX2_51/Y vdd INVX2
XINVX2_73 INVX2_73/A gnd INVX2_73/Y vdd INVX2
XFILL_7_0_0 gnd vdd FILL
XFILL_8_5_1 gnd vdd FILL
XINVX2_62 INVX1_61/A gnd INVX2_62/Y vdd INVX2
XINVX2_40 NOR2X1_1/A gnd OR2X2_1/A vdd INVX2
XINVX2_95 INVX1_36/A gnd INVX2_95/Y vdd INVX2
XFILL_16_4_1 gnd vdd FILL
XINVX2_84 INVX1_55/A gnd INVX2_84/Y vdd INVX2
XOAI21X1_25 INVX1_13/Y BUFX4_161/Y NAND2X1_13/Y gnd NAND3X1_15/B vdd OAI21X1
XOAI21X1_58 BUFX4_183/Y INVX2_13/Y OAI21X1_58/C gnd DFFSR_5/D vdd OAI21X1
XOAI21X1_36 BUFX4_182/Y INVX2_2/Y OAI21X1_36/C gnd DFFSR_10/D vdd OAI21X1
XOAI21X1_69 INVX2_18/Y BUFX4_7/Y OAI21X1_69/C gnd OAI21X1_69/Y vdd OAI21X1
XOAI21X1_14 BUFX4_180/Y INVX1_7/Y NAND3X1_9/Y gnd DFFSR_31/D vdd OAI21X1
XOAI21X1_47 INVX2_8/Y BUFX4_12/Y OAI21X1_47/C gnd NAND3X1_26/B vdd OAI21X1
XOAI21X1_217 NOR2X1_93/Y NOR2X1_94/Y BUFX4_198/Y gnd OAI21X1_217/Y vdd OAI21X1
XOAI21X1_206 NOR2X1_71/Y NOR2X1_72/Y BUFX4_194/Y gnd OAI21X1_206/Y vdd OAI21X1
XOAI21X1_239 NOR2X1_125/Y NOR2X1_126/Y BUFX4_187/Y gnd OAI21X1_239/Y vdd OAI21X1
XOAI21X1_228 DFFSR_172/Q INVX8_10/A OAI21X1_228/C gnd AND2X2_14/A vdd OAI21X1
XNAND2X1_223 INVX1_122/A NOR2X1_189/Y gnd OR2X2_12/B vdd NAND2X1
XNAND2X1_201 wb_dat_i[31] BUFX4_70/Y gnd OAI21X1_738/C vdd NAND2X1
XNAND2X1_212 BUFX4_70/Y wb_dat_i[24] gnd OAI21X1_353/C vdd NAND2X1
XAND2X2_28 AND2X2_28/A INVX4_9/A gnd AND2X2_28/Y vdd AND2X2
XAND2X2_17 NOR2X1_87/B AND2X2_17/B gnd AND2X2_17/Y vdd AND2X2
XNAND2X1_234 INVX1_130/Y INVX8_17/A gnd NAND2X1_234/Y vdd NAND2X1
XNAND2X1_245 BUFX4_81/Y wb_dat_i[1] gnd NAND2X1_245/Y vdd NAND2X1
XNAND2X1_267 INVX2_78/A BUFX4_211/Y gnd NAND2X1_267/Y vdd NAND2X1
XNAND2X1_278 INVX4_10/A NOR2X1_276/Y gnd AOI21X1_234/B vdd NAND2X1
XNAND2X1_289 BUFX4_205/Y NAND2X1_289/B gnd OAI21X1_666/C vdd NAND2X1
XNAND2X1_256 INVX4_8/A AND2X2_23/A gnd NAND2X1_256/Y vdd NAND2X1
XOAI21X1_795 NAND2X1_107/Y INVX4_11/Y OAI21X1_795/C gnd OAI21X1_796/A vdd OAI21X1
XOAI21X1_784 BUFX4_60/Y NAND2X1_338/Y OAI21X1_784/C gnd OAI21X1_784/Y vdd OAI21X1
XOAI21X1_762 BUFX4_220/Y OAI21X1_762/B BUFX4_48/Y gnd AOI21X1_255/A vdd OAI21X1
XOAI21X1_773 INVX2_129/Y BUFX4_164/Y NAND2X1_330/Y gnd AOI21X1_262/B vdd OAI21X1
XOAI21X1_751 AND2X2_31/Y INVX2_126/Y BUFX4_119/Y gnd AOI21X1_252/C vdd OAI21X1
XOAI21X1_740 OAI21X1_740/A OAI21X1_740/B OAI21X1_735/Y gnd DFFSR_211/D vdd OAI21X1
XDFFSR_17 INVX1_9/A DFFSR_2/CLK DFFSR_88/R vdd DFFSR_17/D gnd vdd DFFSR
XFILL_31_2_1 gnd vdd FILL
XDFFSR_28 INVX1_4/A DFFSR_28/CLK DFFSR_25/R vdd DFFSR_28/D gnd vdd DFFSR
XCLKBUF1_15 CLKBUF1_46/A gnd DFFSR_2/CLK vdd CLKBUF1
XDFFSR_39 XOR2X1_3/B CLKBUF1_37/Y DFFSR_2/R vdd DFFSR_39/D gnd vdd DFFSR
XCLKBUF1_37 CLKBUF1_46/A gnd CLKBUF1_37/Y vdd CLKBUF1
XCLKBUF1_48 CLKBUF1_6/A gnd CLKBUF1_48/Y vdd CLKBUF1
XCLKBUF1_59 wb_clk_i gnd CLKBUF1_4/A vdd CLKBUF1
XBUFX4_80 wb_sel_i[0] gnd BUFX4_80/Y vdd BUFX4
XBUFX4_91 INVX8_3/Y gnd BUFX4_91/Y vdd BUFX4
XCLKBUF1_26 CLKBUF1_56/Y gnd CLKBUF1_26/Y vdd CLKBUF1
XFILL_22_2_1 gnd vdd FILL
XXNOR2X1_1 NOR2X1_41/Y XNOR2X1_1/B gnd XNOR2X1_1/Y vdd XNOR2X1
XFILL_5_3_1 gnd vdd FILL
XINVX1_1 INVX1_1/A gnd INVX1_1/Y vdd INVX1
XFILL_13_2_1 gnd vdd FILL
XOAI21X1_592 INVX2_163/Y BUFX4_162/Y NAND2X1_216/Y gnd AOI21X1_202/B vdd OAI21X1
XOAI21X1_581 NOR2X1_273/Y INVX1_138/Y BUFX4_119/Y gnd OAI21X1_581/Y vdd OAI21X1
XOAI21X1_570 BUFX4_96/Y INVX8_11/Y AND2X2_23/A gnd INVX1_139/A vdd OAI21X1
XBUFX4_217 BUFX4_217/A gnd BUFX4_217/Y vdd BUFX4
XBUFX4_206 BUFX4_211/A gnd BUFX4_206/Y vdd BUFX4
XBUFX4_228 BUFX4_228/A gnd OAI22X1_1/D vdd BUFX4
XBUFX4_239 BUFX4_239/A gnd BUFX4_239/Y vdd BUFX4
XAND2X2_1 BUFX4_23/Y AND2X2_1/B gnd AND2X2_1/Y vdd AND2X2
XFILL_2_1 gnd vdd FILL
XNAND3X1_17 BUFX4_19/Y NAND3X1_17/B BUFX4_26/Y gnd OAI21X1_30/C vdd NAND3X1
XNAND3X1_28 BUFX4_16/Y NAND3X1_28/B BUFX4_24/Y gnd NAND3X1_28/Y vdd NAND3X1
XNAND3X1_39 OAI21X1_71/Y BUFX4_18/Y INVX8_2/Y gnd OAI21X1_72/C vdd NAND3X1
XNOR2X1_17 NOR2X1_17/A NOR2X1_17/B gnd NOR2X1_17/Y vdd NOR2X1
XNOR2X1_28 INVX1_72/A DFFSR_107/Q gnd AND2X2_4/A vdd NOR2X1
XFILL_27_1_1 gnd vdd FILL
XFILL_2_1_1 gnd vdd FILL
XNOR2X1_39 XOR2X1_1/A XOR2X1_1/B gnd AND2X2_5/B vdd NOR2X1
XFILL_10_0_1 gnd vdd FILL
XNOR2X1_118 INVX2_107/Y BUFX4_45/Y gnd NOR2X1_118/Y vdd NOR2X1
XNOR2X1_129 INVX2_116/Y NOR2X1_71/B gnd NOR2X1_129/Y vdd NOR2X1
XFILL_18_1_1 gnd vdd FILL
XNOR2X1_107 INVX2_90/Y BUFX4_46/Y gnd NOR2X1_107/Y vdd NOR2X1
XDFFSR_5 DFFSR_5/Q DFFSR_5/CLK DFFSR_1/R vdd DFFSR_5/D gnd vdd DFFSR
XNAND2X1_61 DFFSR_133/Q AOI21X1_1/B gnd NAND3X1_87/A vdd NAND2X1
XNAND2X1_50 NAND3X1_80/Y NAND2X1_50/B gnd AOI21X1_10/C vdd NAND2X1
XNAND2X1_94 INVX1_72/Y AND2X2_5/Y gnd NAND2X1_94/Y vdd NAND2X1
XNAND2X1_72 INVX1_95/A BUFX4_190/Y gnd NAND3X1_98/A vdd NAND2X1
XNAND2X1_83 NOR2X1_1/A BUFX2_2/A gnd NAND2X1_83/Y vdd NAND2X1
XAOI21X1_210 NOR2X1_280/Y BUFX4_61/Y AOI21X1_210/C gnd OAI21X1_601/A vdd AOI21X1
XAOI21X1_232 AOI21X1_231/Y AOI21X1_232/B NOR2X1_289/Y gnd DFFSR_154/D vdd AOI21X1
XAOI21X1_265 INVX2_132/Y OR2X2_21/Y INVX8_15/A gnd OAI21X1_778/C vdd AOI21X1
XAOI21X1_254 INVX2_130/Y NAND2X1_332/Y BUFX4_230/Y gnd OAI21X1_760/C vdd AOI21X1
XAOI21X1_243 MUX2X1_5/B INVX1_142/Y BUFX4_207/Y gnd AOI22X1_78/D vdd AOI21X1
XAOI21X1_221 BUFX4_30/Y AOI21X1_221/B BUFX4_203/Y gnd AOI21X1_222/A vdd AOI21X1
XAOI22X1_81 BUFX4_212/Y MUX2X1_8/Y AOI22X1_81/C AOI22X1_81/D gnd DFFSR_142/D vdd AOI22X1
XAOI22X1_70 INVX2_65/A INVX8_14/A INVX4_8/A INVX2_63/A gnd AOI22X1_70/Y vdd AOI22X1
XNAND3X1_203 OAI21X1_301/Y OAI21X1_302/Y AOI22X1_53/Y gnd AOI22X1_54/C vdd NAND3X1
XDFFSR_212 INVX1_26/A CLKBUF1_13/Y DFFSR_198/R vdd DFFSR_212/D gnd vdd DFFSR
XDFFSR_234 INVX2_52/A CLKBUF1_37/Y DFFSR_198/R vdd DFFSR_234/D gnd vdd DFFSR
XDFFSR_201 INVX2_160/A CLKBUF1_50/Y DFFSR_203/R vdd DFFSR_201/D gnd vdd DFFSR
XDFFSR_223 INVX1_54/A CLKBUF1_24/Y DFFSR_194/R vdd DFFSR_223/D gnd vdd DFFSR
XDFFSR_245 BUFX4_98/A CLKBUF1_4/Y DFFSR_165/R vdd DFFSR_245/D gnd vdd DFFSR
XINVX2_74 INVX2_74/A gnd INVX2_74/Y vdd INVX2
XINVX2_52 INVX2_52/A gnd INVX2_52/Y vdd INVX2
XINVX2_41 INVX2_41/A gnd INVX2_41/Y vdd INVX2
XFILL_7_0_1 gnd vdd FILL
XINVX2_63 INVX2_63/A gnd INVX2_63/Y vdd INVX2
XINVX2_96 INVX2_96/A gnd INVX2_96/Y vdd INVX2
XINVX2_30 INVX2_30/A gnd INVX2_30/Y vdd INVX2
XINVX2_85 INVX1_56/A gnd INVX2_85/Y vdd INVX2
XOAI21X1_26 BUFX4_179/Y INVX1_13/Y OAI21X1_26/C gnd DFFSR_21/D vdd OAI21X1
XOAI21X1_59 INVX2_14/Y BUFX4_82/Y OAI21X1_59/C gnd OAI21X1_59/Y vdd OAI21X1
XOAI21X1_15 INVX1_8/Y MUX2X1_8/S NAND2X1_8/Y gnd NAND3X1_10/B vdd OAI21X1
XOAI21X1_48 BUFX4_182/Y INVX2_8/Y OAI21X1_48/C gnd DFFSR_16/D vdd OAI21X1
XOAI21X1_37 INVX2_3/Y BUFX4_10/Y OAI21X1_67/C gnd NAND3X1_21/B vdd OAI21X1
XAND2X2_18 INVX2_43/A INVX2_48/A gnd AND2X2_18/Y vdd AND2X2
XOAI21X1_218 NOR2X1_95/Y NOR2X1_96/Y BUFX4_198/Y gnd NAND3X1_121/B vdd OAI21X1
XOAI21X1_207 NOR2X1_73/Y NOR2X1_74/Y BUFX4_185/Y gnd OAI21X1_207/Y vdd OAI21X1
XAND2X2_29 AND2X2_29/A INVX4_9/A gnd AND2X2_29/Y vdd AND2X2
XOAI21X1_229 AND2X2_13/Y AND2X2_14/Y NOR2X1_76/B gnd OAI21X1_229/Y vdd OAI21X1
XNAND2X1_268 DFFSR_165/Q BUFX4_204/Y gnd OAI21X1_606/C vdd NAND2X1
XNAND2X1_224 BUFX4_162/Y wb_dat_i[18] gnd NAND2X1_224/Y vdd NAND2X1
XNAND2X1_246 INVX8_17/A INVX1_129/Y gnd AOI21X1_147/B vdd NAND2X1
XNAND2X1_213 INVX1_122/A NOR2X1_190/Y gnd NOR2X1_243/B vdd NAND2X1
XNAND2X1_202 BUFX4_72/Y wb_dat_i[30] gnd OAI21X1_323/C vdd NAND2X1
XNAND2X1_257 INVX2_64/A BUFX4_207/Y gnd NAND2X1_257/Y vdd NAND2X1
XNAND2X1_235 BUFX4_9/Y wb_dat_i[11] gnd OAI21X1_621/C vdd NAND2X1
XNAND2X1_279 INVX4_10/A NOR2X1_278/Y gnd AOI21X1_237/B vdd NAND2X1
XOAI21X1_730 INVX1_160/Y INVX1_99/A BUFX4_113/Y gnd OAI21X1_730/Y vdd OAI21X1
XNOR2X1_290 OR2X2_17/B OR2X2_16/A gnd NOR2X1_290/Y vdd NOR2X1
XOAI21X1_741 BUFX4_222/Y BUFX4_233/Y INVX1_62/A gnd OAI21X1_741/Y vdd OAI21X1
XOAI21X1_796 OAI21X1_796/A INVX4_5/Y NAND2X1_344/Y gnd DFFSR_250/D vdd OAI21X1
XOAI21X1_785 INVX2_131/Y BUFX4_165/Y NAND2X1_330/Y gnd NAND2X1_339/B vdd OAI21X1
XOAI21X1_763 INVX8_21/A BUFX4_28/Y INVX2_134/A gnd OAI21X1_763/Y vdd OAI21X1
XOAI21X1_774 NOR2X1_335/Y INVX2_133/Y BUFX4_120/Y gnd AOI21X1_264/C vdd OAI21X1
XOAI21X1_752 INVX2_126/Y BUFX4_73/Y OAI21X1_738/C gnd OAI21X1_753/B vdd OAI21X1
XDFFSR_18 INVX1_10/A DFFSR_3/CLK DFFSR_7/R vdd DFFSR_18/D gnd vdd DFFSR
XDFFSR_29 INVX1_5/A CLKBUF1_8/A DFFSR_95/R vdd DFFSR_29/D gnd vdd DFFSR
XCLKBUF1_27 CLKBUF1_54/Y gnd CLKBUF1_27/Y vdd CLKBUF1
XCLKBUF1_38 CLKBUF1_38/A gnd DFFSR_99/CLK vdd CLKBUF1
XCLKBUF1_16 CLKBUF1_34/A gnd DFFSR_92/CLK vdd CLKBUF1
XBUFX4_92 INVX8_3/Y gnd BUFX4_92/Y vdd BUFX4
XBUFX4_81 wb_sel_i[0] gnd BUFX4_81/Y vdd BUFX4
XCLKBUF1_49 CLKBUF1_3/A gnd DFFSR_6/CLK vdd CLKBUF1
XBUFX4_70 wb_sel_i[3] gnd BUFX4_70/Y vdd BUFX4
XXNOR2X1_2 NOR2X1_44/B INVX2_41/Y gnd XNOR2X1_2/Y vdd XNOR2X1
XOAI21X1_593 BUFX4_64/Y NAND2X1_265/Y OAI21X1_593/C gnd AOI21X1_206/B vdd OAI21X1
XOAI21X1_560 BUFX4_119/Y OAI21X1_560/B BUFX4_116/Y gnd OAI21X1_561/B vdd OAI21X1
XINVX1_2 INVX1_2/A gnd INVX1_2/Y vdd INVX1
XOAI21X1_571 NOR2X1_271/Y INVX2_68/Y BUFX4_123/Y gnd AOI21X1_197/C vdd OAI21X1
XOAI21X1_582 INVX1_138/Y BUFX4_71/Y OAI21X1_353/C gnd OAI21X1_583/B vdd OAI21X1
XFILL_32_5_0 gnd vdd FILL
XFILL_23_5_0 gnd vdd FILL
XBUFX4_207 BUFX4_211/A gnd BUFX4_207/Y vdd BUFX4
XFILL_6_6_0 gnd vdd FILL
XBUFX4_218 BUFX4_217/A gnd NOR2X1_87/B vdd BUFX4
XBUFX4_229 BUFX4_230/A gnd BUFX4_229/Y vdd BUFX4
XFILL_14_5_0 gnd vdd FILL
XAND2X2_2 INVX8_2/Y AND2X2_2/B gnd AND2X2_2/Y vdd AND2X2
XOAI21X1_390 NOR2X1_220/Y INVX2_84/Y BUFX4_54/Y gnd OAI21X1_390/Y vdd OAI21X1
XFILL_2_2 gnd vdd FILL
XNAND3X1_18 BUFX4_19/Y NAND3X1_18/B BUFX4_24/Y gnd NAND3X1_18/Y vdd NAND3X1
XNOR2X1_18 BUFX2_35/A NOR2X1_18/B gnd DFFSR_64/D vdd NOR2X1
XNAND3X1_29 BUFX4_15/Y OAI21X1_53/Y BUFX4_24/Y gnd NAND3X1_29/Y vdd NAND3X1
XNOR2X1_29 XNOR2X1_1/B DFFSR_106/Q gnd AND2X2_4/B vdd NOR2X1
XNOR2X1_108 INVX2_91/Y BUFX4_215/Y gnd NOR2X1_108/Y vdd NOR2X1
XNOR2X1_119 INVX2_108/Y NOR2X1_99/B gnd NOR2X1_119/Y vdd NOR2X1
XDFFSR_6 DFFSR_6/Q DFFSR_6/CLK DFFSR_7/R vdd DFFSR_6/D gnd vdd DFFSR
XNAND2X1_62 INVX2_80/A AOI21X1_1/B gnd NAND2X1_62/Y vdd NAND2X1
XNAND2X1_40 NAND3X1_73/Y NAND2X1_40/B gnd AOI21X1_3/C vdd NAND2X1
XNAND2X1_51 NAND2X1_51/A NOR2X1_13/Y gnd DFFSR_74/D vdd NAND2X1
XNAND2X1_73 MUX2X1_5/B BUFX4_192/Y gnd NAND3X1_99/B vdd NAND2X1
XNAND2X1_95 INVX2_37/A BUFX4_3/Y gnd NAND2X1_95/Y vdd NAND2X1
XNAND2X1_84 AND2X2_5/A AND2X2_5/B gnd NOR3X1_2/C vdd NAND2X1
XAOI21X1_200 NOR2X1_274/Y BUFX4_58/Y AOI21X1_200/C gnd OAI21X1_589/A vdd AOI21X1
XAOI21X1_211 NOR2X1_281/Y BUFX4_58/Y AOI21X1_211/C gnd OAI21X1_606/A vdd AOI21X1
XAOI21X1_233 NOR2X1_290/Y BUFX4_58/Y AOI21X1_233/C gnd OAI21X1_635/A vdd AOI21X1
XAOI21X1_266 BUFX4_150/Y AOI21X1_266/B BUFX4_48/Y gnd AOI21X1_267/A vdd AOI21X1
XFILL_20_3_0 gnd vdd FILL
XAOI21X1_255 AOI21X1_255/A AOI21X1_255/B NOR2X1_331/Y gnd DFFSR_203/D vdd AOI21X1
XAOI21X1_244 INVX1_95/A INVX1_143/Y BUFX4_212/Y gnd AOI22X1_79/D vdd AOI21X1
XAOI22X1_82 BUFX4_212/Y MUX2X1_9/Y AOI22X1_82/C AOI22X1_82/D gnd DFFSR_127/D vdd AOI22X1
XAOI22X1_60 INVX2_126/A INVX4_9/A INVX8_23/A INVX1_98/A gnd AOI22X1_60/Y vdd AOI22X1
XAOI22X1_71 INVX2_61/A INVX4_10/A INVX8_22/A INVX1_92/A gnd AOI22X1_71/Y vdd AOI22X1
XAOI21X1_222 AOI21X1_222/A AOI21X1_222/B NOR2X1_285/Y gnd DFFSR_159/D vdd AOI21X1
XFILL_28_4_0 gnd vdd FILL
XFILL_3_4_0 gnd vdd FILL
XNAND3X1_204 OAI21X1_304/Y NAND3X1_204/B AOI22X1_55/Y gnd AOI22X1_57/A vdd NAND3X1
XFILL_11_3_0 gnd vdd FILL
XFILL_19_4_0 gnd vdd FILL
XDFFSR_246 OR2X2_8/A DFFSR_36/CLK BUFX4_130/Y vdd DFFSR_246/D gnd vdd DFFSR
XDFFSR_202 INVX2_55/A CLKBUF1_48/Y BUFX4_130/Y vdd DFFSR_202/D gnd vdd DFFSR
XDFFSR_213 INVX1_28/A CLKBUF1_11/Y DFFSR_198/R vdd DFFSR_213/D gnd vdd DFFSR
XDFFSR_224 INVX1_55/A CLKBUF1_56/Y DFFSR_236/R vdd DFFSR_224/D gnd vdd DFFSR
XDFFSR_235 INVX2_128/A CLKBUF1_33/Y DFFSR_203/R vdd DFFSR_235/D gnd vdd DFFSR
XINVX2_42 INVX2_42/A gnd INVX2_42/Y vdd INVX2
XINVX2_53 XOR2X1_3/A gnd INVX2_53/Y vdd INVX2
XINVX2_20 INVX2_49/A gnd INVX2_20/Y vdd INVX2
XINVX2_75 INVX1_30/A gnd INVX2_75/Y vdd INVX2
XINVX2_31 OR2X2_2/B gnd INVX2_31/Y vdd INVX2
XINVX2_64 INVX2_64/A gnd INVX2_64/Y vdd INVX2
XINVX2_86 INVX2_86/A gnd INVX2_86/Y vdd INVX2
XINVX2_97 INVX1_47/A gnd INVX2_97/Y vdd INVX2
XOAI21X1_16 BUFX4_182/Y INVX1_8/Y OAI21X1_16/C gnd DFFSR_32/D vdd OAI21X1
XOAI21X1_27 INVX1_14/Y BUFX4_163/Y OAI21X1_27/C gnd NAND3X1_16/B vdd OAI21X1
XOAI21X1_49 INVX2_9/Y BUFX4_80/Y NAND2X1_25/Y gnd OAI21X1_49/Y vdd OAI21X1
XOAI21X1_38 BUFX4_182/Y INVX2_3/Y OAI21X1_38/C gnd DFFSR_11/D vdd OAI21X1
XFILL_34_2_0 gnd vdd FILL
XOAI21X1_219 NOR2X1_97/Y NOR2X1_98/Y BUFX4_184/Y gnd NAND3X1_121/C vdd OAI21X1
XOAI21X1_208 NOR2X1_76/Y NOR2X1_75/Y AND2X2_16/B gnd OAI21X1_208/Y vdd OAI21X1
XAND2X2_19 INVX2_42/A INVX8_13/A gnd AND2X2_19/Y vdd AND2X2
XNAND2X1_269 DFFSR_164/Q BUFX4_204/Y gnd NAND2X1_269/Y vdd NAND2X1
XNAND2X1_214 wb_dat_i[22] BUFX4_161/Y gnd OAI21X1_587/C vdd NAND2X1
XNAND2X1_247 BUFX4_83/Y wb_dat_i[0] gnd OAI21X1_732/C vdd NAND2X1
XNAND2X1_225 INVX1_125/Y NOR2X1_189/Y gnd OR2X2_13/B vdd NAND2X1
XNAND2X1_203 MUX2X1_6/S wb_dat_i[29] gnd OAI21X1_328/C vdd NAND2X1
XNAND2X1_258 INVX4_9/A NOR2X1_266/Y gnd NAND2X1_258/Y vdd NAND2X1
XNAND2X1_236 BUFX4_11/Y wb_dat_i[10] gnd NAND2X1_236/Y vdd NAND2X1
XFILL_25_2_0 gnd vdd FILL
XFILL_0_2_0 gnd vdd FILL
XOAI21X1_731 NOR2X1_323/Y OAI21X1_730/Y NAND2X1_324/Y gnd DFFSR_117/D vdd OAI21X1
XNOR2X1_280 INVX4_9/Y NOR2X1_280/B gnd NOR2X1_280/Y vdd NOR2X1
XOAI21X1_775 INVX2_133/Y BUFX4_84/Y OAI21X1_787/C gnd OAI21X1_776/B vdd OAI21X1
XOAI21X1_764 AND2X2_32/Y INVX2_134/Y BUFX4_169/Y gnd OAI21X1_764/Y vdd OAI21X1
XNOR2X1_291 INVX1_35/A BUFX4_115/Y gnd NOR2X1_291/Y vdd NOR2X1
XOAI21X1_720 BUFX4_60/Y NAND2X1_319/Y OAI21X1_720/C gnd OAI21X1_720/Y vdd OAI21X1
XOAI21X1_753 BUFX4_123/Y OAI21X1_753/B BUFX4_116/Y gnd OAI21X1_754/B vdd OAI21X1
XOAI21X1_742 NOR2X1_326/Y INVX2_122/Y BUFX4_56/Y gnd AOI21X1_250/C vdd OAI21X1
XOAI21X1_797 OR2X2_7/B INVX4_11/A BUFX4_101/Y gnd OAI22X1_45/D vdd OAI21X1
XOAI21X1_786 OAI21X1_784/Y BUFX4_206/Y OAI21X1_786/C gnd DFFSR_139/D vdd OAI21X1
XFILL_8_3_0 gnd vdd FILL
XFILL_16_2_0 gnd vdd FILL
XDFFSR_19 INVX1_11/A CLKBUF1_5/Y DFFSR_1/R vdd DFFSR_19/D gnd vdd DFFSR
XCLKBUF1_28 CLKBUF1_34/A gnd CLKBUF1_28/Y vdd CLKBUF1
XCLKBUF1_17 CLKBUF1_5/A gnd DFFSR_46/CLK vdd CLKBUF1
XCLKBUF1_39 CLKBUF1_5/A gnd CLKBUF1_39/Y vdd CLKBUF1
XBUFX4_93 INVX8_3/Y gnd BUFX4_93/Y vdd BUFX4
XBUFX4_82 wb_sel_i[0] gnd BUFX4_82/Y vdd BUFX4
XBUFX4_60 BUFX4_61/A gnd BUFX4_60/Y vdd BUFX4
XBUFX4_71 wb_sel_i[3] gnd BUFX4_71/Y vdd BUFX4
XXNOR2X1_3 OR2X2_8/B INVX2_46/A gnd XNOR2X1_3/Y vdd XNOR2X1
XOR2X2_1 OR2X2_1/A BUFX2_2/A gnd OR2X2_1/Y vdd OR2X2
XOAI21X1_550 INVX2_146/Y BUFX4_82/Y NAND2X1_245/Y gnd OAI21X1_551/B vdd OAI21X1
XOAI21X1_594 INVX2_88/Y BUFX4_163/Y NAND2X1_219/Y gnd AOI21X1_205/B vdd OAI21X1
XINVX1_3 INVX1_3/A gnd INVX1_3/Y vdd INVX1
XOAI21X1_561 OAI21X1_561/A OAI21X1_561/B NAND2X1_257/Y gnd DFFSR_178/D vdd OAI21X1
XOAI21X1_572 INVX2_68/Y MUX2X1_8/S OAI21X1_572/C gnd OAI21X1_573/B vdd OAI21X1
XOAI21X1_583 BUFX4_123/Y OAI21X1_583/B BUFX4_116/Y gnd OAI21X1_583/Y vdd OAI21X1
XFILL_32_5_1 gnd vdd FILL
XFILL_31_0_0 gnd vdd FILL
XFILL_23_5_1 gnd vdd FILL
XFILL_22_0_0 gnd vdd FILL
XBUFX4_208 BUFX4_211/A gnd BUFX4_208/Y vdd BUFX4
XBUFX4_219 BUFX4_217/A gnd NOR2X1_71/B vdd BUFX4
XFILL_5_1_0 gnd vdd FILL
XFILL_6_6_1 gnd vdd FILL
XFILL_13_0_0 gnd vdd FILL
XFILL_14_5_1 gnd vdd FILL
XOAI21X1_380 BUFX4_66/Y AOI21X1_121/B OAI21X1_380/C gnd OAI21X1_380/Y vdd OAI21X1
XAND2X2_3 AND2X2_3/A BUFX4_20/Y gnd AND2X2_3/Y vdd AND2X2
XOAI21X1_391 INVX2_84/Y BUFX4_8/Y OAI21X1_699/C gnd OAI21X1_392/B vdd OAI21X1
XNAND3X1_19 BUFX4_18/Y OAI21X1_33/Y BUFX4_27/Y gnd OAI21X1_34/C vdd NAND3X1
XNOR2X1_19 NOR2X1_1/B NOR2X1_19/B gnd NOR2X1_19/Y vdd NOR2X1
XNOR2X1_109 INVX2_92/Y BUFX4_42/Y gnd NOR2X1_109/Y vdd NOR2X1
XDFFSR_7 DFFSR_7/Q DFFSR_7/CLK DFFSR_7/R vdd DFFSR_7/D gnd vdd DFFSR
XNAND2X1_30 BUFX4_81/Y wb_dat_i[5] gnd OAI21X1_59/C vdd NAND2X1
XNAND2X1_41 AOI21X1_3/Y NOR2X1_6/Y gnd DFFSR_67/D vdd NAND2X1
XNAND2X1_63 DFFSR_135/Q AOI21X1_7/B gnd NAND2X1_63/Y vdd NAND2X1
XNAND2X1_52 NAND2X1_52/A NAND2X1_52/B gnd AOI21X1_11/C vdd NAND2X1
XNAND2X1_74 INVX1_92/A BUFX4_192/Y gnd NAND2X1_74/Y vdd NAND2X1
XNAND2X1_96 DFFSR_54/Q BUFX4_3/Y gnd NAND2X1_96/Y vdd NAND2X1
XNAND2X1_85 BUFX2_2/A NAND2X1_85/B gnd NAND2X1_85/Y vdd NAND2X1
XAOI21X1_212 NOR2X1_282/Y BUFX4_61/Y AOI21X1_212/C gnd AOI21X1_212/Y vdd AOI21X1
XAOI21X1_201 INVX2_163/Y OR2X2_16/Y BUFX4_32/Y gnd OAI21X1_591/C vdd AOI21X1
XFILL_20_3_1 gnd vdd FILL
XAOI21X1_234 INVX2_92/Y AOI21X1_234/B BUFX4_33/Y gnd OAI21X1_636/C vdd AOI21X1
XAOI21X1_223 INVX2_71/Y AOI21X1_223/B BUFX4_34/Y gnd OAI21X1_622/C vdd AOI21X1
XAOI21X1_256 AND2X2_32/Y BUFX4_66/Y OAI21X1_764/Y gnd AOI21X1_256/Y vdd AOI21X1
XAOI21X1_267 AOI21X1_267/A AOI21X1_267/B NOR2X1_336/Y gnd DFFSR_219/D vdd AOI21X1
XAOI22X1_50 NOR2X1_189/Y AOI22X1_50/B AOI22X1_50/C INVX2_164/A gnd AOI21X1_85/A vdd
+ AOI22X1
XAOI21X1_245 INVX1_96/A INVX1_144/Y BUFX4_212/Y gnd AOI22X1_80/D vdd AOI21X1
XAOI22X1_83 BUFX4_210/Y MUX2X1_10/Y AOI22X1_83/C AOI22X1_83/D gnd DFFSR_126/D vdd
+ AOI22X1
XAOI22X1_61 DFFSR_163/Q INVX4_10/A INVX4_8/A INVX1_63/A gnd AOI22X1_61/Y vdd AOI22X1
XAOI22X1_72 INVX1_61/A INVX8_17/A INVX8_23/A INVX1_91/A gnd AOI22X1_72/Y vdd AOI22X1
XFILL_28_4_1 gnd vdd FILL
XNAND3X1_205 NAND3X1_205/A NAND3X1_205/B AOI22X1_56/Y gnd AOI22X1_57/D vdd NAND3X1
XFILL_3_4_1 gnd vdd FILL
XFILL_11_3_1 gnd vdd FILL
XOAI22X1_1 BUFX4_78/Y INVX2_9/Y INVX1_26/Y OAI22X1_1/D gnd NOR2X1_2/A vdd OAI22X1
XFILL_19_4_1 gnd vdd FILL
XDFFSR_247 OR2X2_8/B CLKBUF1_48/Y BUFX4_130/Y vdd DFFSR_247/D gnd vdd DFFSR
XDFFSR_214 INVX1_30/A CLKBUF1_6/Y BUFX4_130/Y vdd DFFSR_214/D gnd vdd DFFSR
XDFFSR_203 INVX2_130/A CLKBUF1_42/Y DFFSR_203/R vdd DFFSR_203/D gnd vdd DFFSR
XDFFSR_225 INVX1_59/A CLKBUF1_32/A DFFSR_236/R vdd DFFSR_225/D gnd vdd DFFSR
XDFFSR_236 INVX2_165/A CLKBUF1_32/Y DFFSR_236/R vdd DFFSR_236/D gnd vdd DFFSR
XINVX2_10 DFFSR_2/Q gnd INVX2_10/Y vdd INVX2
XINVX2_21 INVX2_50/A gnd INVX2_21/Y vdd INVX2
XINVX2_43 INVX2_43/A gnd INVX2_43/Y vdd INVX2
XINVX2_54 INVX2_54/A gnd INVX2_54/Y vdd INVX2
XINVX2_76 INVX1_31/A gnd INVX2_76/Y vdd INVX2
XINVX2_32 INVX2_32/A gnd INVX2_32/Y vdd INVX2
XINVX2_87 INVX2_87/A gnd INVX2_87/Y vdd INVX2
XINVX2_65 INVX2_65/A gnd INVX2_65/Y vdd INVX2
XINVX2_98 INVX2_98/A gnd INVX2_98/Y vdd INVX2
XOAI21X1_17 INVX1_9/Y BUFX4_160/Y NAND2X1_9/Y gnd NAND3X1_11/B vdd OAI21X1
XOAI21X1_28 BUFX4_179/Y INVX1_14/Y OAI21X1_28/C gnd DFFSR_22/D vdd OAI21X1
XOAI21X1_39 INVX2_4/Y BUFX4_12/Y OAI21X1_69/C gnd OAI21X1_39/Y vdd OAI21X1
XFILL_34_2_1 gnd vdd FILL
XOAI21X1_209 NOR2X1_78/Y NOR2X1_77/Y BUFX4_188/Y gnd OAI21X1_209/Y vdd OAI21X1
XNAND2X1_226 BUFX4_164/Y wb_dat_i[17] gnd NAND2X1_226/Y vdd NAND2X1
XNAND2X1_215 INVX1_125/Y NOR2X1_190/Y gnd NOR2X1_245/B vdd NAND2X1
XNAND2X1_204 MUX2X1_8/S wb_dat_i[28] gnd OAI21X1_333/C vdd NAND2X1
XNAND2X1_248 INVX4_7/A INVX1_131/Y gnd NAND2X1_248/Y vdd NAND2X1
XNAND2X1_259 INVX4_9/A AND2X2_30/A gnd NAND2X1_259/Y vdd NAND2X1
XNAND2X1_237 BUFX4_5/Y wb_dat_i[9] gnd OAI21X1_515/C vdd NAND2X1
XNOR2X1_281 INVX4_9/Y NOR2X1_310/B gnd NOR2X1_281/Y vdd NOR2X1
XNOR2X1_292 INVX1_32/A BUFX4_114/Y gnd NOR2X1_292/Y vdd NOR2X1
XFILL_25_2_1 gnd vdd FILL
XFILL_0_2_1 gnd vdd FILL
XNOR2X1_270 BUFX4_229/Y INVX1_133/A gnd AND2X2_29/A vdd NOR2X1
XOAI21X1_798 OR2X2_7/Y INVX4_11/Y XOR2X1_3/A gnd AOI21X1_268/A vdd OAI21X1
XOAI21X1_732 INVX2_107/Y BUFX4_81/Y OAI21X1_732/C gnd OAI21X1_732/Y vdd OAI21X1
XOAI21X1_787 INVX2_135/Y BUFX4_86/Y OAI21X1_787/C gnd OAI21X1_787/Y vdd OAI21X1
XOAI21X1_765 INVX2_134/Y BUFX4_83/Y OAI21X1_787/C gnd OAI21X1_765/Y vdd OAI21X1
XOAI21X1_776 BUFX4_120/Y OAI21X1_776/B BUFX4_115/Y gnd OAI21X1_777/B vdd OAI21X1
XOAI21X1_721 OAI21X1_720/Y BUFX4_208/Y NAND2X1_318/Y gnd DFFSR_120/D vdd OAI21X1
XOAI21X1_754 OAI21X1_754/A OAI21X1_754/B NAND2X1_331/Y gnd DFFSR_179/D vdd OAI21X1
XOAI21X1_710 OAI21X1_710/A BUFX4_210/Y OAI21X1_710/C gnd DFFSR_124/D vdd OAI21X1
XOAI21X1_743 INVX2_122/Y BUFX4_7/Y NAND2X1_328/Y gnd OAI21X1_744/B vdd OAI21X1
XFILL_8_3_1 gnd vdd FILL
XFILL_16_2_1 gnd vdd FILL
XCLKBUF1_29 CLKBUF1_4/A gnd DFFSR_71/CLK vdd CLKBUF1
XCLKBUF1_18 CLKBUF1_3/A gnd DFFSR_1/CLK vdd CLKBUF1
XBUFX4_61 BUFX4_61/A gnd BUFX4_61/Y vdd BUFX4
XBUFX4_50 BUFX4_47/A gnd BUFX4_50/Y vdd BUFX4
XBUFX4_83 wb_sel_i[0] gnd BUFX4_83/Y vdd BUFX4
XBUFX4_94 INVX8_3/Y gnd BUFX4_94/Y vdd BUFX4
XBUFX4_72 wb_sel_i[3] gnd BUFX4_72/Y vdd BUFX4
XXNOR2X1_4 INVX2_43/A INVX4_2/A gnd XNOR2X1_4/Y vdd XNOR2X1
XOR2X2_20 OR2X2_20/A INVX4_9/Y gnd OR2X2_20/Y vdd OR2X2
XOR2X2_2 OR2X2_2/A OR2X2_2/B gnd OR2X2_2/Y vdd OR2X2
XINVX8_20 BUFX4_32/Y gnd INVX8_20/Y vdd INVX8
XINVX1_4 INVX1_4/A gnd INVX1_4/Y vdd INVX1
XOAI21X1_551 BUFX4_170/Y OAI21X1_551/B BUFX4_36/Y gnd OAI21X1_552/B vdd OAI21X1
XOAI21X1_540 INVX2_116/Y BUFX4_80/Y NAND2X1_243/Y gnd OAI21X1_540/Y vdd OAI21X1
XOAI21X1_595 BUFX4_64/Y NAND2X1_266/Y OAI21X1_595/C gnd AOI21X1_209/B vdd OAI21X1
XOAI21X1_562 BUFX4_63/Y NAND2X1_258/Y AOI21X1_190/Y gnd OAI21X1_562/Y vdd OAI21X1
XOAI21X1_573 BUFX4_123/Y OAI21X1_573/B BUFX4_117/Y gnd OAI21X1_574/B vdd OAI21X1
XOAI21X1_584 OAI21X1_584/A OAI21X1_583/Y NAND2X1_263/Y gnd DFFSR_172/D vdd OAI21X1
XFILL_31_0_1 gnd vdd FILL
XFILL_22_0_1 gnd vdd FILL
XBUFX4_209 BUFX4_211/A gnd INVX8_21/A vdd BUFX4
XFILL_5_1_1 gnd vdd FILL
XFILL_13_0_1 gnd vdd FILL
XOAI21X1_381 INVX2_102/Y BUFX4_160/Y NAND2X1_229/Y gnd OAI21X1_381/Y vdd OAI21X1
XOAI21X1_370 BUFX4_221/Y BUFX4_230/Y INVX2_77/A gnd OAI21X1_374/C vdd OAI21X1
XAND2X2_4 AND2X2_4/A AND2X2_4/B gnd AND2X2_4/Y vdd AND2X2
XOAI21X1_392 BUFX4_54/Y OAI21X1_392/B BUFX4_242/Y gnd OAI21X1_392/Y vdd OAI21X1
XDFFSR_8 DFFSR_8/Q DFFSR_8/CLK DFFSR_9/R vdd DFFSR_8/D gnd vdd DFFSR
XNAND2X1_31 BUFX4_83/Y wb_dat_i[6] gnd OAI21X1_90/C vdd NAND2X1
XNAND2X1_64 INVX2_90/A AOI21X1_2/B gnd NAND2X1_64/Y vdd NAND2X1
XNAND2X1_42 AOI21X1_4/Y NOR2X1_7/Y gnd DFFSR_68/D vdd NAND2X1
XNAND2X1_75 AND2X2_17/B BUFX4_192/Y gnd NAND2X1_75/Y vdd NAND2X1
XNAND2X1_86 AND2X2_4/Y AND2X2_5/Y gnd NAND2X1_86/Y vdd NAND2X1
XNAND2X1_97 INVX2_24/A BUFX4_2/Y gnd NAND2X1_97/Y vdd NAND2X1
XNAND2X1_53 NAND2X1_53/A NOR2X1_14/Y gnd DFFSR_75/D vdd NAND2X1
XNAND2X1_20 BUFX4_11/Y wb_dat_i[11] gnd OAI21X1_69/C vdd NAND2X1
XAOI21X1_202 BUFX4_32/Y AOI21X1_202/B BUFX4_206/Y gnd AOI21X1_202/Y vdd AOI21X1
XAOI21X1_235 BUFX4_33/Y OAI21X1_637/Y BUFX4_208/Y gnd AOI21X1_235/Y vdd AOI21X1
XAOI21X1_257 AND2X2_17/B INVX1_162/Y BUFX4_212/Y gnd AOI22X1_84/D vdd AOI21X1
XAOI21X1_246 INVX1_93/A INVX1_145/Y BUFX4_212/Y gnd AOI22X1_81/D vdd AOI21X1
XAOI21X1_224 BUFX4_34/Y AOI21X1_224/B BUFX4_205/Y gnd AOI21X1_225/A vdd AOI21X1
XAOI21X1_213 INVX2_61/Y NAND2X1_270/Y BUFX4_30/Y gnd OAI21X1_612/C vdd AOI21X1
XAOI21X1_268 AOI21X1_268/A NOR2X1_346/Y AND2X2_33/A gnd DFFSR_252/D vdd AOI21X1
XAOI22X1_51 AOI22X1_51/A AOI21X1_77/Y AOI22X1_51/C AOI22X1_51/D gnd AOI22X1_51/Y vdd
+ AOI22X1
XAOI22X1_84 BUFX4_212/Y MUX2X1_11/Y AOI22X1_84/C AOI22X1_84/D gnd DFFSR_147/D vdd
+ AOI22X1
XAOI22X1_62 INVX2_109/A INVX4_9/A INVX4_7/A INVX2_110/A gnd AOI22X1_62/Y vdd AOI22X1
XAOI22X1_73 INVX1_50/A INVX8_17/A INVX4_7/A INVX2_69/A gnd AOI22X1_73/Y vdd AOI22X1
XAOI22X1_40 AOI22X1_40/A AOI21X1_58/Y AOI22X1_40/C AOI22X1_40/D gnd AOI22X1_40/Y vdd
+ AOI22X1
XNAND3X1_206 OAI21X1_308/Y OAI21X1_309/Y AOI22X1_57/Y gnd AOI22X1_77/A vdd NAND3X1
XOAI22X1_2 OAI22X1_4/A INVX2_31/Y OAI22X1_4/C INVX1_27/Y gnd NOR2X1_2/B vdd OAI22X1
XFILL_30_6_0 gnd vdd FILL
XDFFSR_248 INVX2_43/A DFFSR_83/CLK BUFX4_130/Y vdd DFFSR_248/D gnd vdd DFFSR
XDFFSR_215 INVX1_34/A CLKBUF1_1/Y DFFSR_203/R vdd DFFSR_215/D gnd vdd DFFSR
XDFFSR_237 INVX2_141/A CLKBUF1_26/Y DFFSR_236/R vdd DFFSR_237/D gnd vdd DFFSR
XDFFSR_204 DFFSR_204/Q CLKBUF1_39/Y DFFSR_167/R vdd DFFSR_204/D gnd vdd DFFSR
XDFFSR_226 INVX1_61/A CLKBUF1_19/Y DFFSR_203/R vdd DFFSR_226/D gnd vdd DFFSR
XFILL_21_6_0 gnd vdd FILL
XINVX2_11 DFFSR_3/Q gnd INVX2_11/Y vdd INVX2
XINVX2_22 XOR2X1_3/B gnd INVX2_22/Y vdd INVX2
XINVX2_44 OR2X2_8/A gnd INVX2_44/Y vdd INVX2
XINVX2_33 INVX2_33/A gnd INVX2_33/Y vdd INVX2
XINVX2_55 INVX2_55/A gnd INVX2_55/Y vdd INVX2
XINVX2_77 INVX2_77/A gnd INVX2_77/Y vdd INVX2
XINVX2_88 INVX2_88/A gnd INVX2_88/Y vdd INVX2
XINVX2_66 INVX2_66/A gnd INVX2_66/Y vdd INVX2
XINVX2_99 INVX1_46/A gnd INVX2_99/Y vdd INVX2
XOAI21X1_18 BUFX4_179/Y INVX1_9/Y OAI21X1_18/C gnd DFFSR_17/D vdd OAI21X1
XOAI21X1_29 INVX1_15/Y BUFX4_165/Y OAI21X1_29/C gnd NAND3X1_17/B vdd OAI21X1
XFILL_12_6_0 gnd vdd FILL
XNAND2X1_216 BUFX4_163/Y wb_dat_i[21] gnd NAND2X1_216/Y vdd NAND2X1
XNAND2X1_205 INVX1_111/A NOR2X1_191/Y gnd INVX1_130/A vdd NAND2X1
XNAND2X1_227 INVX1_126/Y NOR2X1_189/Y gnd INVX1_129/A vdd NAND2X1
XNAND2X1_238 BUFX4_7/Y wb_dat_i[8] gnd NAND2X1_238/Y vdd NAND2X1
XNAND2X1_249 INVX4_7/A INVX1_133/Y gnd NAND2X1_249/Y vdd NAND2X1
XNOR2X1_282 INVX4_9/Y NOR2X1_282/B gnd NOR2X1_282/Y vdd NOR2X1
XNOR2X1_293 OR2X2_17/B NOR2X1_280/B gnd NOR2X1_293/Y vdd NOR2X1
XNOR2X1_271 INVX4_9/Y INVX1_139/A gnd NOR2X1_271/Y vdd NOR2X1
XNOR2X1_260 INVX4_8/Y INVX1_134/Y gnd NOR2X1_260/Y vdd NOR2X1
XOAI21X1_799 AOI22X1_85/C NAND2X1_345/Y AOI22X1_85/Y gnd DFFSR_253/D vdd OAI21X1
XOAI21X1_733 INVX1_161/Y DFFSR_116/Q BUFX4_113/Y gnd OAI21X1_733/Y vdd OAI21X1
XOAI21X1_766 BUFX4_170/Y OAI21X1_765/Y BUFX4_37/Y gnd OAI21X1_766/Y vdd OAI21X1
XOAI21X1_711 INVX1_149/Y OR2X2_18/B INVX2_60/Y gnd OAI21X1_711/Y vdd OAI21X1
XOAI21X1_777 OAI21X1_777/A OAI21X1_777/B NAND2X1_336/Y gnd DFFSR_155/D vdd OAI21X1
XOAI21X1_788 INVX1_164/Y OR2X2_18/B INVX2_135/Y gnd OAI21X1_788/Y vdd OAI21X1
XOAI21X1_722 INVX2_117/Y BUFX4_86/Y NAND2X1_243/Y gnd NAND2X1_320/B vdd OAI21X1
XOAI21X1_700 OR2X2_18/A OR2X2_18/B INVX2_87/Y gnd OAI21X1_700/Y vdd OAI21X1
XOAI21X1_744 BUFX4_56/Y OAI21X1_744/B BUFX4_240/Y gnd OAI21X1_744/Y vdd OAI21X1
XOAI21X1_755 BUFX4_205/Y BUFX4_29/Y INVX1_63/A gnd OAI21X1_755/Y vdd OAI21X1
XBUFX4_95 INVX8_3/Y gnd BUFX4_95/Y vdd BUFX4
XBUFX4_84 wb_sel_i[0] gnd BUFX4_84/Y vdd BUFX4
XCLKBUF1_19 CLKBUF1_5/A gnd CLKBUF1_19/Y vdd CLKBUF1
XBUFX4_73 wb_sel_i[3] gnd BUFX4_73/Y vdd BUFX4
XBUFX4_62 BUFX4_61/A gnd BUFX4_62/Y vdd BUFX4
XBUFX4_40 BUFX4_45/A gnd BUFX4_40/Y vdd BUFX4
XBUFX4_51 BUFX4_52/A gnd BUFX4_51/Y vdd BUFX4
XFILL_35_5_0 gnd vdd FILL
XOR2X2_10 OR2X2_10/A DFFSR_33/Q gnd OR2X2_10/Y vdd OR2X2
XOR2X2_21 OR2X2_12/A OR2X2_21/B gnd OR2X2_21/Y vdd OR2X2
XXNOR2X1_5 OR2X2_7/Y INVX2_53/Y gnd INVX1_89/A vdd XNOR2X1
XOR2X2_3 BUFX2_2/A OR2X2_3/B gnd OR2X2_3/Y vdd OR2X2
XFILL_26_5_0 gnd vdd FILL
XFILL_1_5_0 gnd vdd FILL
XOAI21X1_541 BUFX4_169/Y OAI21X1_540/Y BUFX4_37/Y gnd OAI21X1_541/Y vdd OAI21X1
XOAI21X1_530 INVX2_157/Y BUFX4_86/Y NAND2X1_240/Y gnd OAI21X1_531/B vdd OAI21X1
XINVX8_21 INVX8_21/A gnd INVX8_21/Y vdd INVX8
XINVX8_10 INVX8_10/A gnd INVX8_10/Y vdd INVX8
XINVX1_5 INVX1_5/A gnd INVX1_5/Y vdd INVX1
XOAI21X1_552 AOI21X1_187/Y OAI21X1_552/B OAI21X1_552/C gnd DFFSR_181/D vdd OAI21X1
XOAI21X1_585 BUFX4_98/Y INVX8_11/Y AND2X2_25/A gnd OR2X2_17/A vdd OAI21X1
XOAI21X1_596 INVX2_121/Y BUFX4_164/Y NAND2X1_222/Y gnd OAI21X1_596/Y vdd OAI21X1
XOAI21X1_563 INVX2_151/Y BUFX4_73/Y OAI21X1_328/C gnd AOI21X1_191/B vdd OAI21X1
XOAI21X1_574 OAI21X1_574/A OAI21X1_574/B NAND2X1_261/Y gnd DFFSR_174/D vdd OAI21X1
.ends

